library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"c248d4ff",
     1 => x"78bff1f5",
     2 => x"bfedf5c2",
     3 => x"edf5c249",
     4 => x"78a1c148",
     5 => x"a9b7c0c4",
     6 => x"ff87e504",
     7 => x"78c848d0",
     8 => x"48f9f5c2",
     9 => x"4f2678c0",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"5f000000",
    13 => x"0000005f",
    14 => x"00030300",
    15 => x"00000303",
    16 => x"147f7f14",
    17 => x"00147f7f",
    18 => x"6b2e2400",
    19 => x"00123a6b",
    20 => x"18366a4c",
    21 => x"0032566c",
    22 => x"594f7e30",
    23 => x"40683a77",
    24 => x"07040000",
    25 => x"00000003",
    26 => x"3e1c0000",
    27 => x"00004163",
    28 => x"63410000",
    29 => x"00001c3e",
    30 => x"1c3e2a08",
    31 => x"082a3e1c",
    32 => x"3e080800",
    33 => x"0008083e",
    34 => x"e0800000",
    35 => x"00000060",
    36 => x"08080800",
    37 => x"00080808",
    38 => x"60000000",
    39 => x"00000060",
    40 => x"18306040",
    41 => x"0103060c",
    42 => x"597f3e00",
    43 => x"003e7f4d",
    44 => x"7f060400",
    45 => x"0000007f",
    46 => x"71634200",
    47 => x"00464f59",
    48 => x"49632200",
    49 => x"00367f49",
    50 => x"13161c18",
    51 => x"00107f7f",
    52 => x"45672700",
    53 => x"00397d45",
    54 => x"4b7e3c00",
    55 => x"00307949",
    56 => x"71010100",
    57 => x"00070f79",
    58 => x"497f3600",
    59 => x"00367f49",
    60 => x"494f0600",
    61 => x"001e3f69",
    62 => x"66000000",
    63 => x"00000066",
    64 => x"e6800000",
    65 => x"00000066",
    66 => x"14080800",
    67 => x"00222214",
    68 => x"14141400",
    69 => x"00141414",
    70 => x"14222200",
    71 => x"00080814",
    72 => x"51030200",
    73 => x"00060f59",
    74 => x"5d417f3e",
    75 => x"001e1f55",
    76 => x"097f7e00",
    77 => x"007e7f09",
    78 => x"497f7f00",
    79 => x"00367f49",
    80 => x"633e1c00",
    81 => x"00414141",
    82 => x"417f7f00",
    83 => x"001c3e63",
    84 => x"497f7f00",
    85 => x"00414149",
    86 => x"097f7f00",
    87 => x"00010109",
    88 => x"417f3e00",
    89 => x"007a7b49",
    90 => x"087f7f00",
    91 => x"007f7f08",
    92 => x"7f410000",
    93 => x"0000417f",
    94 => x"40602000",
    95 => x"003f7f40",
    96 => x"1c087f7f",
    97 => x"00416336",
    98 => x"407f7f00",
    99 => x"00404040",
   100 => x"0c067f7f",
   101 => x"007f7f06",
   102 => x"0c067f7f",
   103 => x"007f7f18",
   104 => x"417f3e00",
   105 => x"003e7f41",
   106 => x"097f7f00",
   107 => x"00060f09",
   108 => x"61417f3e",
   109 => x"00407e7f",
   110 => x"097f7f00",
   111 => x"00667f19",
   112 => x"4d6f2600",
   113 => x"00327b59",
   114 => x"7f010100",
   115 => x"0001017f",
   116 => x"407f3f00",
   117 => x"003f7f40",
   118 => x"703f0f00",
   119 => x"000f3f70",
   120 => x"18307f7f",
   121 => x"007f7f30",
   122 => x"1c366341",
   123 => x"4163361c",
   124 => x"7c060301",
   125 => x"0103067c",
   126 => x"4d597161",
   127 => x"00414347",
   128 => x"7f7f0000",
   129 => x"00004141",
   130 => x"0c060301",
   131 => x"40603018",
   132 => x"41410000",
   133 => x"00007f7f",
   134 => x"03060c08",
   135 => x"00080c06",
   136 => x"80808080",
   137 => x"00808080",
   138 => x"03000000",
   139 => x"00000407",
   140 => x"54742000",
   141 => x"00787c54",
   142 => x"447f7f00",
   143 => x"00387c44",
   144 => x"447c3800",
   145 => x"00004444",
   146 => x"447c3800",
   147 => x"007f7f44",
   148 => x"547c3800",
   149 => x"00185c54",
   150 => x"7f7e0400",
   151 => x"00000505",
   152 => x"a4bc1800",
   153 => x"007cfca4",
   154 => x"047f7f00",
   155 => x"00787c04",
   156 => x"3d000000",
   157 => x"0000407d",
   158 => x"80808000",
   159 => x"00007dfd",
   160 => x"107f7f00",
   161 => x"00446c38",
   162 => x"3f000000",
   163 => x"0000407f",
   164 => x"180c7c7c",
   165 => x"00787c0c",
   166 => x"047c7c00",
   167 => x"00787c04",
   168 => x"447c3800",
   169 => x"00387c44",
   170 => x"24fcfc00",
   171 => x"00183c24",
   172 => x"243c1800",
   173 => x"00fcfc24",
   174 => x"047c7c00",
   175 => x"00080c04",
   176 => x"545c4800",
   177 => x"00207454",
   178 => x"7f3f0400",
   179 => x"00004444",
   180 => x"407c3c00",
   181 => x"007c7c40",
   182 => x"603c1c00",
   183 => x"001c3c60",
   184 => x"30607c3c",
   185 => x"003c7c60",
   186 => x"10386c44",
   187 => x"00446c38",
   188 => x"e0bc1c00",
   189 => x"001c3c60",
   190 => x"74644400",
   191 => x"00444c5c",
   192 => x"3e080800",
   193 => x"00414177",
   194 => x"7f000000",
   195 => x"0000007f",
   196 => x"77414100",
   197 => x"0008083e",
   198 => x"03010102",
   199 => x"00010202",
   200 => x"7f7f7f7f",
   201 => x"007f7f7f",
   202 => x"1c1c0808",
   203 => x"7f7f3e3e",
   204 => x"3e3e7f7f",
   205 => x"08081c1c",
   206 => x"7c181000",
   207 => x"0010187c",
   208 => x"7c301000",
   209 => x"0010307c",
   210 => x"60603010",
   211 => x"00061e78",
   212 => x"183c6642",
   213 => x"0042663c",
   214 => x"c26a3878",
   215 => x"00386cc6",
   216 => x"60000060",
   217 => x"00600000",
   218 => x"5c5b5e0e",
   219 => x"711e0e5d",
   220 => x"caf6c24c",
   221 => x"4bc04dbf",
   222 => x"ab741ec0",
   223 => x"c487c702",
   224 => x"78c048a6",
   225 => x"a6c487c5",
   226 => x"c478c148",
   227 => x"49731e66",
   228 => x"c887dfee",
   229 => x"49e0c086",
   230 => x"c487efef",
   231 => x"496a4aa5",
   232 => x"f187f0f0",
   233 => x"85cb87c6",
   234 => x"b7c883c1",
   235 => x"c7ff04ab",
   236 => x"4d262687",
   237 => x"4b264c26",
   238 => x"711e4f26",
   239 => x"cef6c24a",
   240 => x"cef6c25a",
   241 => x"4978c748",
   242 => x"2687ddfe",
   243 => x"1e731e4f",
   244 => x"b7c04a71",
   245 => x"87d303aa",
   246 => x"bfeddcc2",
   247 => x"c187c405",
   248 => x"c087c24b",
   249 => x"f1dcc24b",
   250 => x"c287c45b",
   251 => x"c25af1dc",
   252 => x"4abfeddc",
   253 => x"c0c19ac1",
   254 => x"e8ec49a2",
   255 => x"c248fc87",
   256 => x"78bfeddc",
   257 => x"1e87effe",
   258 => x"66c44a71",
   259 => x"ff49721e",
   260 => x"2687dadf",
   261 => x"c21e4f26",
   262 => x"49bfeddc",
   263 => x"87c2dcff",
   264 => x"48c2f6c2",
   265 => x"c278bfe8",
   266 => x"ec48fef5",
   267 => x"f6c278bf",
   268 => x"494abfc2",
   269 => x"c899ffc3",
   270 => x"48722ab7",
   271 => x"f6c2b071",
   272 => x"4f2658ca",
   273 => x"5c5b5e0e",
   274 => x"4b710e5d",
   275 => x"c287c7ff",
   276 => x"c048fdf5",
   277 => x"ff497350",
   278 => x"7087e7db",
   279 => x"9cc24c49",
   280 => x"cb49eecb",
   281 => x"497087cf",
   282 => x"fdf5c24d",
   283 => x"c105bf97",
   284 => x"66d087e4",
   285 => x"c6f6c249",
   286 => x"d70599bf",
   287 => x"4966d487",
   288 => x"bffef5c2",
   289 => x"87cc0599",
   290 => x"daff4973",
   291 => x"987087f4",
   292 => x"87c2c102",
   293 => x"fdfd4cc1",
   294 => x"ca497587",
   295 => x"987087e3",
   296 => x"c287c602",
   297 => x"c148fdf5",
   298 => x"fdf5c250",
   299 => x"c005bf97",
   300 => x"f6c287e4",
   301 => x"d049bfc6",
   302 => x"ff059966",
   303 => x"f5c287d6",
   304 => x"d449bffe",
   305 => x"ff059966",
   306 => x"497387ca",
   307 => x"87f2d9ff",
   308 => x"fe059870",
   309 => x"487487fe",
   310 => x"0e87d7fb",
   311 => x"5d5c5b5e",
   312 => x"c086f40e",
   313 => x"bfec4c4d",
   314 => x"48a6c47e",
   315 => x"bfcaf6c2",
   316 => x"c01ec178",
   317 => x"fd49c71e",
   318 => x"86c887ca",
   319 => x"ce029870",
   320 => x"fb49ff87",
   321 => x"dac187c7",
   322 => x"f5d8ff49",
   323 => x"c24dc187",
   324 => x"bf97fdf5",
   325 => x"cd87c302",
   326 => x"f6c287f9",
   327 => x"c24bbfc2",
   328 => x"05bfeddc",
   329 => x"c387ebc0",
   330 => x"d8ff49fd",
   331 => x"fac387d4",
   332 => x"cdd8ff49",
   333 => x"c3497387",
   334 => x"1e7199ff",
   335 => x"c6fb49c0",
   336 => x"c8497387",
   337 => x"1e7129b7",
   338 => x"fafa49c1",
   339 => x"c686c887",
   340 => x"f6c287c1",
   341 => x"9b4bbfc6",
   342 => x"c287dd02",
   343 => x"49bfe9dc",
   344 => x"7087dec7",
   345 => x"87c40598",
   346 => x"87d24bc0",
   347 => x"c749e0c2",
   348 => x"dcc287c3",
   349 => x"87c658ed",
   350 => x"48e9dcc2",
   351 => x"497378c0",
   352 => x"ce0599c2",
   353 => x"49ebc387",
   354 => x"87f6d6ff",
   355 => x"99c24970",
   356 => x"fb87c202",
   357 => x"c149734c",
   358 => x"87ce0599",
   359 => x"ff49f4c3",
   360 => x"7087dfd6",
   361 => x"0299c249",
   362 => x"4cfa87c2",
   363 => x"99c84973",
   364 => x"c387ce05",
   365 => x"d6ff49f5",
   366 => x"497087c8",
   367 => x"d50299c2",
   368 => x"cef6c287",
   369 => x"87ca02bf",
   370 => x"c288c148",
   371 => x"c058d2f6",
   372 => x"4cff87c2",
   373 => x"49734dc1",
   374 => x"ce0599c4",
   375 => x"49f2c387",
   376 => x"87ded5ff",
   377 => x"99c24970",
   378 => x"c287dc02",
   379 => x"7ebfcef6",
   380 => x"a8b7c748",
   381 => x"87cbc003",
   382 => x"80c1486e",
   383 => x"58d2f6c2",
   384 => x"fe87c2c0",
   385 => x"c34dc14c",
   386 => x"d4ff49fd",
   387 => x"497087f4",
   388 => x"c00299c2",
   389 => x"f6c287d5",
   390 => x"c002bfce",
   391 => x"f6c287c9",
   392 => x"78c048ce",
   393 => x"fd87c2c0",
   394 => x"c34dc14c",
   395 => x"d4ff49fa",
   396 => x"497087d0",
   397 => x"c00299c2",
   398 => x"f6c287d9",
   399 => x"c748bfce",
   400 => x"c003a8b7",
   401 => x"f6c287c9",
   402 => x"78c748ce",
   403 => x"fc87c2c0",
   404 => x"c04dc14c",
   405 => x"c003acb7",
   406 => x"66c487d1",
   407 => x"82d8c14a",
   408 => x"c6c0026a",
   409 => x"744b6a87",
   410 => x"c00f7349",
   411 => x"1ef0c31e",
   412 => x"f749dac1",
   413 => x"86c887ce",
   414 => x"c0029870",
   415 => x"a6c887e2",
   416 => x"cef6c248",
   417 => x"66c878bf",
   418 => x"c491cb49",
   419 => x"80714866",
   420 => x"bf6e7e70",
   421 => x"87c8c002",
   422 => x"c84bbf6e",
   423 => x"0f734966",
   424 => x"c0029d75",
   425 => x"f6c287c8",
   426 => x"f249bfce",
   427 => x"dcc287fa",
   428 => x"c002bff1",
   429 => x"c24987dd",
   430 => x"987087c7",
   431 => x"87d3c002",
   432 => x"bfcef6c2",
   433 => x"87e0f249",
   434 => x"c0f449c0",
   435 => x"f1dcc287",
   436 => x"f478c048",
   437 => x"87daf38e",
   438 => x"5c5b5e0e",
   439 => x"711e0e5d",
   440 => x"caf6c24c",
   441 => x"cdc149bf",
   442 => x"d1c14da1",
   443 => x"747e6981",
   444 => x"87cf029c",
   445 => x"744ba5c4",
   446 => x"caf6c27b",
   447 => x"f9f249bf",
   448 => x"747b6e87",
   449 => x"87c4059c",
   450 => x"87c24bc0",
   451 => x"49734bc1",
   452 => x"d487faf2",
   453 => x"87c70266",
   454 => x"7087da49",
   455 => x"c087c24a",
   456 => x"f5dcc24a",
   457 => x"c9f2265a",
   458 => x"00000087",
   459 => x"00000000",
   460 => x"00000000",
   461 => x"4a711e00",
   462 => x"49bfc8ff",
   463 => x"2648a172",
   464 => x"c8ff1e4f",
   465 => x"c0fe89bf",
   466 => x"c0c0c0c0",
   467 => x"87c401a9",
   468 => x"87c24ac0",
   469 => x"48724ac1",
   470 => x"5e0e4f26",
   471 => x"0e5d5c5b",
   472 => x"ff4d711e",
   473 => x"1e754bd4",
   474 => x"49d2f6c2",
   475 => x"87f2c1fe",
   476 => x"7e7086c4",
   477 => x"ffc3026e",
   478 => x"daf6c287",
   479 => x"49754cbf",
   480 => x"87e0dbfe",
   481 => x"c005a8de",
   482 => x"497587eb",
   483 => x"87ecd3ff",
   484 => x"db029870",
   485 => x"d5f5c287",
   486 => x"e1c01ebf",
   487 => x"f7d0ff49",
   488 => x"c286c487",
   489 => x"c048d2e2",
   490 => x"e1f5c250",
   491 => x"87eafe49",
   492 => x"c5c348c1",
   493 => x"48d0ff87",
   494 => x"c178c5c8",
   495 => x"4ac07bd6",
   496 => x"7bbf976e",
   497 => x"80c1486e",
   498 => x"82c17e70",
   499 => x"aab7e0c0",
   500 => x"87ecff04",
   501 => x"c448d0ff",
   502 => x"78c5c878",
   503 => x"c17bd3c1",
   504 => x"7478c47b",
   505 => x"fdc1029c",
   506 => x"cee4c287",
   507 => x"4dc0c87e",
   508 => x"acb7c08c",
   509 => x"c887c603",
   510 => x"c04da4c0",
   511 => x"fff0c24c",
   512 => x"d049bf97",
   513 => x"87d20299",
   514 => x"f6c21ec0",
   515 => x"c2fe49d2",
   516 => x"86c487ec",
   517 => x"c04a4970",
   518 => x"e4c287ef",
   519 => x"f6c21ece",
   520 => x"c2fe49d2",
   521 => x"86c487d8",
   522 => x"ff4a4970",
   523 => x"c5c848d0",
   524 => x"7bd4c178",
   525 => x"7bbf976e",
   526 => x"80c1486e",
   527 => x"8dc17e70",
   528 => x"87f0ff05",
   529 => x"c448d0ff",
   530 => x"059a7278",
   531 => x"c087c5c0",
   532 => x"87e6c048",
   533 => x"f6c21ec1",
   534 => x"fffd49d2",
   535 => x"86c487ff",
   536 => x"fe059c74",
   537 => x"d0ff87c3",
   538 => x"78c5c848",
   539 => x"c07bd3c1",
   540 => x"c178c47b",
   541 => x"87c2c048",
   542 => x"262648c0",
   543 => x"264c264d",
   544 => x"1e4f264b",
   545 => x"66c44a71",
   546 => x"7287c505",
   547 => x"87cafb49",
   548 => x"1e004f26",
   549 => x"bfe1e3c2",
   550 => x"c2b9c149",
   551 => x"ff59e5e3",
   552 => x"ffc348d4",
   553 => x"48d0ff78",
   554 => x"ff78e1c8",
   555 => x"78c148d4",
   556 => x"787131c4",
   557 => x"c048d0ff",
   558 => x"4f2678e0",
   559 => x"d5e3c21e",
   560 => x"d2f6c21e",
   561 => x"d9fcfd49",
   562 => x"7086c487",
   563 => x"87c30298",
   564 => x"2687c0ff",
   565 => x"4b35314f",
   566 => x"20205a48",
   567 => x"47464320",
   568 => x"00000000",
   569 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
