
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"f6",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"e8",x"f6",x"c2"),
    14 => (x"48",x"e8",x"e3",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ff",x"df"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"ff",x"1e",x"4f",x"26"),
    53 => (x"ff",x"c3",x"48",x"d4"),
    54 => (x"c4",x"51",x"68",x"78"),
    55 => (x"88",x"c1",x"48",x"66"),
    56 => (x"70",x"58",x"a6",x"c8"),
    57 => (x"87",x"eb",x"05",x"98"),
    58 => (x"73",x"1e",x"4f",x"26"),
    59 => (x"4b",x"d4",x"ff",x"1e"),
    60 => (x"6b",x"7b",x"ff",x"c3"),
    61 => (x"7b",x"ff",x"c3",x"4a"),
    62 => (x"32",x"c8",x"49",x"6b"),
    63 => (x"ff",x"c3",x"b1",x"72"),
    64 => (x"c8",x"4a",x"6b",x"7b"),
    65 => (x"c3",x"b2",x"71",x"31"),
    66 => (x"49",x"6b",x"7b",x"ff"),
    67 => (x"b1",x"72",x"32",x"c8"),
    68 => (x"87",x"c4",x"48",x"71"),
    69 => (x"4c",x"26",x"4d",x"26"),
    70 => (x"4f",x"26",x"4b",x"26"),
    71 => (x"5c",x"5b",x"5e",x"0e"),
    72 => (x"4a",x"71",x"0e",x"5d"),
    73 => (x"72",x"4c",x"d4",x"ff"),
    74 => (x"99",x"ff",x"c3",x"49"),
    75 => (x"e3",x"c2",x"7c",x"71"),
    76 => (x"c8",x"05",x"bf",x"e8"),
    77 => (x"48",x"66",x"d0",x"87"),
    78 => (x"a6",x"d4",x"30",x"c9"),
    79 => (x"49",x"66",x"d0",x"58"),
    80 => (x"ff",x"c3",x"29",x"d8"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"d0",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"ff",x"c3",x"29",x"c8"),
    86 => (x"d0",x"7c",x"71",x"99"),
    87 => (x"ff",x"c3",x"49",x"66"),
    88 => (x"72",x"7c",x"71",x"99"),
    89 => (x"c3",x"29",x"d0",x"49"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"f0",x"c9",x"4b",x"6c"),
    92 => (x"ff",x"c3",x"4d",x"ff"),
    93 => (x"87",x"d0",x"05",x"ab"),
    94 => (x"6c",x"7c",x"ff",x"c3"),
    95 => (x"02",x"8d",x"c1",x"4b"),
    96 => (x"ff",x"c3",x"87",x"c6"),
    97 => (x"87",x"f0",x"02",x"ab"),
    98 => (x"c7",x"fe",x"48",x"73"),
    99 => (x"49",x"c0",x"1e",x"87"),
   100 => (x"c3",x"48",x"d4",x"ff"),
   101 => (x"81",x"c1",x"78",x"ff"),
   102 => (x"a9",x"b7",x"c8",x"c3"),
   103 => (x"26",x"87",x"f1",x"04"),
   104 => (x"1e",x"73",x"1e",x"4f"),
   105 => (x"f8",x"c4",x"87",x"e7"),
   106 => (x"1e",x"c0",x"4b",x"df"),
   107 => (x"c1",x"f0",x"ff",x"c0"),
   108 => (x"e7",x"fd",x"49",x"f7"),
   109 => (x"c1",x"86",x"c4",x"87"),
   110 => (x"ea",x"c0",x"05",x"a8"),
   111 => (x"48",x"d4",x"ff",x"87"),
   112 => (x"c1",x"78",x"ff",x"c3"),
   113 => (x"c0",x"c0",x"c0",x"c0"),
   114 => (x"e1",x"c0",x"1e",x"c0"),
   115 => (x"49",x"e9",x"c1",x"f0"),
   116 => (x"c4",x"87",x"c9",x"fd"),
   117 => (x"05",x"98",x"70",x"86"),
   118 => (x"d4",x"ff",x"87",x"ca"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"87",x"cb",x"48",x"c1"),
   121 => (x"c1",x"87",x"e6",x"fe"),
   122 => (x"fd",x"fe",x"05",x"8b"),
   123 => (x"fc",x"48",x"c0",x"87"),
   124 => (x"73",x"1e",x"87",x"e6"),
   125 => (x"48",x"d4",x"ff",x"1e"),
   126 => (x"d3",x"78",x"ff",x"c3"),
   127 => (x"c0",x"1e",x"c0",x"4b"),
   128 => (x"c1",x"c1",x"f0",x"ff"),
   129 => (x"87",x"d4",x"fc",x"49"),
   130 => (x"98",x"70",x"86",x"c4"),
   131 => (x"ff",x"87",x"ca",x"05"),
   132 => (x"ff",x"c3",x"48",x"d4"),
   133 => (x"cb",x"48",x"c1",x"78"),
   134 => (x"87",x"f1",x"fd",x"87"),
   135 => (x"ff",x"05",x"8b",x"c1"),
   136 => (x"48",x"c0",x"87",x"db"),
   137 => (x"0e",x"87",x"f1",x"fb"),
   138 => (x"0e",x"5c",x"5b",x"5e"),
   139 => (x"fd",x"4c",x"d4",x"ff"),
   140 => (x"ea",x"c6",x"87",x"db"),
   141 => (x"f0",x"e1",x"c0",x"1e"),
   142 => (x"fb",x"49",x"c8",x"c1"),
   143 => (x"86",x"c4",x"87",x"de"),
   144 => (x"c8",x"02",x"a8",x"c1"),
   145 => (x"87",x"ea",x"fe",x"87"),
   146 => (x"e2",x"c1",x"48",x"c0"),
   147 => (x"87",x"da",x"fa",x"87"),
   148 => (x"ff",x"cf",x"49",x"70"),
   149 => (x"ea",x"c6",x"99",x"ff"),
   150 => (x"87",x"c8",x"02",x"a9"),
   151 => (x"c0",x"87",x"d3",x"fe"),
   152 => (x"87",x"cb",x"c1",x"48"),
   153 => (x"c0",x"7c",x"ff",x"c3"),
   154 => (x"f4",x"fc",x"4b",x"f1"),
   155 => (x"02",x"98",x"70",x"87"),
   156 => (x"c0",x"87",x"eb",x"c0"),
   157 => (x"f0",x"ff",x"c0",x"1e"),
   158 => (x"fa",x"49",x"fa",x"c1"),
   159 => (x"86",x"c4",x"87",x"de"),
   160 => (x"d9",x"05",x"98",x"70"),
   161 => (x"7c",x"ff",x"c3",x"87"),
   162 => (x"ff",x"c3",x"49",x"6c"),
   163 => (x"7c",x"7c",x"7c",x"7c"),
   164 => (x"02",x"99",x"c0",x"c1"),
   165 => (x"48",x"c1",x"87",x"c4"),
   166 => (x"48",x"c0",x"87",x"d5"),
   167 => (x"ab",x"c2",x"87",x"d1"),
   168 => (x"c0",x"87",x"c4",x"05"),
   169 => (x"c1",x"87",x"c8",x"48"),
   170 => (x"fd",x"fe",x"05",x"8b"),
   171 => (x"f9",x"48",x"c0",x"87"),
   172 => (x"73",x"1e",x"87",x"e4"),
   173 => (x"e8",x"e3",x"c2",x"1e"),
   174 => (x"c7",x"78",x"c1",x"48"),
   175 => (x"48",x"d0",x"ff",x"4b"),
   176 => (x"c8",x"fb",x"78",x"c2"),
   177 => (x"48",x"d0",x"ff",x"87"),
   178 => (x"1e",x"c0",x"78",x"c3"),
   179 => (x"c1",x"d0",x"e5",x"c0"),
   180 => (x"c7",x"f9",x"49",x"c0"),
   181 => (x"c1",x"86",x"c4",x"87"),
   182 => (x"87",x"c1",x"05",x"a8"),
   183 => (x"05",x"ab",x"c2",x"4b"),
   184 => (x"48",x"c0",x"87",x"c5"),
   185 => (x"c1",x"87",x"f9",x"c0"),
   186 => (x"d0",x"ff",x"05",x"8b"),
   187 => (x"87",x"f7",x"fc",x"87"),
   188 => (x"58",x"ec",x"e3",x"c2"),
   189 => (x"cd",x"05",x"98",x"70"),
   190 => (x"c0",x"1e",x"c1",x"87"),
   191 => (x"d0",x"c1",x"f0",x"ff"),
   192 => (x"87",x"d8",x"f8",x"49"),
   193 => (x"d4",x"ff",x"86",x"c4"),
   194 => (x"78",x"ff",x"c3",x"48"),
   195 => (x"c2",x"87",x"fe",x"c2"),
   196 => (x"ff",x"58",x"f0",x"e3"),
   197 => (x"78",x"c2",x"48",x"d0"),
   198 => (x"c3",x"48",x"d4",x"ff"),
   199 => (x"48",x"c1",x"78",x"ff"),
   200 => (x"1e",x"87",x"f5",x"f7"),
   201 => (x"ff",x"4a",x"d4",x"ff"),
   202 => (x"d1",x"c4",x"48",x"d0"),
   203 => (x"7a",x"ff",x"c3",x"78"),
   204 => (x"f8",x"05",x"89",x"c1"),
   205 => (x"1e",x"4f",x"26",x"87"),
   206 => (x"4b",x"71",x"1e",x"73"),
   207 => (x"df",x"cd",x"ee",x"c5"),
   208 => (x"48",x"d4",x"ff",x"4a"),
   209 => (x"68",x"78",x"ff",x"c3"),
   210 => (x"a8",x"fe",x"c3",x"48"),
   211 => (x"c1",x"87",x"c5",x"02"),
   212 => (x"87",x"ed",x"05",x"8a"),
   213 => (x"c5",x"05",x"9a",x"72"),
   214 => (x"c0",x"48",x"c0",x"87"),
   215 => (x"9b",x"73",x"87",x"ea"),
   216 => (x"c8",x"87",x"cc",x"02"),
   217 => (x"49",x"73",x"1e",x"66"),
   218 => (x"c4",x"87",x"e7",x"f5"),
   219 => (x"c8",x"87",x"c6",x"86"),
   220 => (x"ee",x"fe",x"49",x"66"),
   221 => (x"48",x"d4",x"ff",x"87"),
   222 => (x"78",x"78",x"ff",x"c3"),
   223 => (x"c5",x"05",x"9b",x"73"),
   224 => (x"48",x"d0",x"ff",x"87"),
   225 => (x"48",x"c1",x"78",x"d0"),
   226 => (x"1e",x"87",x"cd",x"f6"),
   227 => (x"4a",x"71",x"1e",x"73"),
   228 => (x"d4",x"ff",x"4b",x"c0"),
   229 => (x"78",x"ff",x"c3",x"48"),
   230 => (x"c4",x"48",x"d0",x"ff"),
   231 => (x"d4",x"ff",x"78",x"c3"),
   232 => (x"78",x"ff",x"c3",x"48"),
   233 => (x"ff",x"c0",x"1e",x"72"),
   234 => (x"49",x"d1",x"c1",x"f0"),
   235 => (x"c4",x"87",x"ed",x"f5"),
   236 => (x"05",x"98",x"70",x"86"),
   237 => (x"c0",x"c8",x"87",x"cd"),
   238 => (x"49",x"66",x"cc",x"1e"),
   239 => (x"c4",x"87",x"f8",x"fd"),
   240 => (x"ff",x"4b",x"70",x"86"),
   241 => (x"78",x"c2",x"48",x"d0"),
   242 => (x"cb",x"f5",x"48",x"73"),
   243 => (x"5b",x"5e",x"0e",x"87"),
   244 => (x"c0",x"0e",x"5d",x"5c"),
   245 => (x"f0",x"ff",x"c0",x"1e"),
   246 => (x"f4",x"49",x"c9",x"c1"),
   247 => (x"1e",x"d2",x"87",x"fe"),
   248 => (x"49",x"f0",x"e3",x"c2"),
   249 => (x"c8",x"87",x"d0",x"fd"),
   250 => (x"c1",x"4c",x"c0",x"86"),
   251 => (x"ac",x"b7",x"d2",x"84"),
   252 => (x"c2",x"87",x"f8",x"04"),
   253 => (x"bf",x"97",x"f0",x"e3"),
   254 => (x"99",x"c0",x"c3",x"49"),
   255 => (x"05",x"a9",x"c0",x"c1"),
   256 => (x"c2",x"87",x"e7",x"c0"),
   257 => (x"bf",x"97",x"f7",x"e3"),
   258 => (x"c2",x"31",x"d0",x"49"),
   259 => (x"bf",x"97",x"f8",x"e3"),
   260 => (x"72",x"32",x"c8",x"4a"),
   261 => (x"f9",x"e3",x"c2",x"b1"),
   262 => (x"b1",x"4a",x"bf",x"97"),
   263 => (x"ff",x"cf",x"4c",x"71"),
   264 => (x"c1",x"9c",x"ff",x"ff"),
   265 => (x"c1",x"34",x"ca",x"84"),
   266 => (x"e3",x"c2",x"87",x"e7"),
   267 => (x"49",x"bf",x"97",x"f9"),
   268 => (x"99",x"c6",x"31",x"c1"),
   269 => (x"97",x"fa",x"e3",x"c2"),
   270 => (x"b7",x"c7",x"4a",x"bf"),
   271 => (x"c2",x"b1",x"72",x"2a"),
   272 => (x"bf",x"97",x"f5",x"e3"),
   273 => (x"9d",x"cf",x"4d",x"4a"),
   274 => (x"97",x"f6",x"e3",x"c2"),
   275 => (x"9a",x"c3",x"4a",x"bf"),
   276 => (x"e3",x"c2",x"32",x"ca"),
   277 => (x"4b",x"bf",x"97",x"f7"),
   278 => (x"b2",x"73",x"33",x"c2"),
   279 => (x"97",x"f8",x"e3",x"c2"),
   280 => (x"c0",x"c3",x"4b",x"bf"),
   281 => (x"2b",x"b7",x"c6",x"9b"),
   282 => (x"81",x"c2",x"b2",x"73"),
   283 => (x"30",x"71",x"48",x"c1"),
   284 => (x"48",x"c1",x"49",x"70"),
   285 => (x"4d",x"70",x"30",x"75"),
   286 => (x"84",x"c1",x"4c",x"72"),
   287 => (x"c0",x"c8",x"94",x"71"),
   288 => (x"cc",x"06",x"ad",x"b7"),
   289 => (x"b7",x"34",x"c1",x"87"),
   290 => (x"b7",x"c0",x"c8",x"2d"),
   291 => (x"f4",x"ff",x"01",x"ad"),
   292 => (x"f1",x"48",x"74",x"87"),
   293 => (x"5e",x"0e",x"87",x"fe"),
   294 => (x"0e",x"5d",x"5c",x"5b"),
   295 => (x"ec",x"c2",x"86",x"f8"),
   296 => (x"78",x"c0",x"48",x"d6"),
   297 => (x"1e",x"ce",x"e4",x"c2"),
   298 => (x"de",x"fb",x"49",x"c0"),
   299 => (x"70",x"86",x"c4",x"87"),
   300 => (x"87",x"c5",x"05",x"98"),
   301 => (x"ce",x"c9",x"48",x"c0"),
   302 => (x"c1",x"4d",x"c0",x"87"),
   303 => (x"ca",x"f5",x"c0",x"7e"),
   304 => (x"e5",x"c2",x"49",x"bf"),
   305 => (x"c8",x"71",x"4a",x"c4"),
   306 => (x"87",x"de",x"ee",x"4b"),
   307 => (x"c2",x"05",x"98",x"70"),
   308 => (x"c0",x"7e",x"c0",x"87"),
   309 => (x"49",x"bf",x"c6",x"f5"),
   310 => (x"4a",x"e0",x"e5",x"c2"),
   311 => (x"ee",x"4b",x"c8",x"71"),
   312 => (x"98",x"70",x"87",x"c8"),
   313 => (x"c0",x"87",x"c2",x"05"),
   314 => (x"c0",x"02",x"6e",x"7e"),
   315 => (x"eb",x"c2",x"87",x"fd"),
   316 => (x"c2",x"4d",x"bf",x"d4"),
   317 => (x"bf",x"9f",x"cc",x"ec"),
   318 => (x"d6",x"c5",x"48",x"7e"),
   319 => (x"c7",x"05",x"a8",x"ea"),
   320 => (x"d4",x"eb",x"c2",x"87"),
   321 => (x"87",x"ce",x"4d",x"bf"),
   322 => (x"e9",x"ca",x"48",x"6e"),
   323 => (x"c5",x"02",x"a8",x"d5"),
   324 => (x"c7",x"48",x"c0",x"87"),
   325 => (x"e4",x"c2",x"87",x"f1"),
   326 => (x"49",x"75",x"1e",x"ce"),
   327 => (x"c4",x"87",x"ec",x"f9"),
   328 => (x"05",x"98",x"70",x"86"),
   329 => (x"48",x"c0",x"87",x"c5"),
   330 => (x"c0",x"87",x"dc",x"c7"),
   331 => (x"49",x"bf",x"c6",x"f5"),
   332 => (x"4a",x"e0",x"e5",x"c2"),
   333 => (x"ec",x"4b",x"c8",x"71"),
   334 => (x"98",x"70",x"87",x"f0"),
   335 => (x"c2",x"87",x"c8",x"05"),
   336 => (x"c1",x"48",x"d6",x"ec"),
   337 => (x"c0",x"87",x"da",x"78"),
   338 => (x"49",x"bf",x"ca",x"f5"),
   339 => (x"4a",x"c4",x"e5",x"c2"),
   340 => (x"ec",x"4b",x"c8",x"71"),
   341 => (x"98",x"70",x"87",x"d4"),
   342 => (x"87",x"c5",x"c0",x"02"),
   343 => (x"e6",x"c6",x"48",x"c0"),
   344 => (x"cc",x"ec",x"c2",x"87"),
   345 => (x"c1",x"49",x"bf",x"97"),
   346 => (x"c0",x"05",x"a9",x"d5"),
   347 => (x"ec",x"c2",x"87",x"cd"),
   348 => (x"49",x"bf",x"97",x"cd"),
   349 => (x"02",x"a9",x"ea",x"c2"),
   350 => (x"c0",x"87",x"c5",x"c0"),
   351 => (x"87",x"c7",x"c6",x"48"),
   352 => (x"97",x"ce",x"e4",x"c2"),
   353 => (x"c3",x"48",x"7e",x"bf"),
   354 => (x"c0",x"02",x"a8",x"e9"),
   355 => (x"48",x"6e",x"87",x"ce"),
   356 => (x"02",x"a8",x"eb",x"c3"),
   357 => (x"c0",x"87",x"c5",x"c0"),
   358 => (x"87",x"eb",x"c5",x"48"),
   359 => (x"97",x"d9",x"e4",x"c2"),
   360 => (x"05",x"99",x"49",x"bf"),
   361 => (x"c2",x"87",x"cc",x"c0"),
   362 => (x"bf",x"97",x"da",x"e4"),
   363 => (x"02",x"a9",x"c2",x"49"),
   364 => (x"c0",x"87",x"c5",x"c0"),
   365 => (x"87",x"cf",x"c5",x"48"),
   366 => (x"97",x"db",x"e4",x"c2"),
   367 => (x"ec",x"c2",x"48",x"bf"),
   368 => (x"4c",x"70",x"58",x"d2"),
   369 => (x"c2",x"88",x"c1",x"48"),
   370 => (x"c2",x"58",x"d6",x"ec"),
   371 => (x"bf",x"97",x"dc",x"e4"),
   372 => (x"c2",x"81",x"75",x"49"),
   373 => (x"bf",x"97",x"dd",x"e4"),
   374 => (x"72",x"32",x"c8",x"4a"),
   375 => (x"f0",x"c2",x"7e",x"a1"),
   376 => (x"78",x"6e",x"48",x"e3"),
   377 => (x"97",x"de",x"e4",x"c2"),
   378 => (x"a6",x"c8",x"48",x"bf"),
   379 => (x"d6",x"ec",x"c2",x"58"),
   380 => (x"d4",x"c2",x"02",x"bf"),
   381 => (x"c6",x"f5",x"c0",x"87"),
   382 => (x"e5",x"c2",x"49",x"bf"),
   383 => (x"c8",x"71",x"4a",x"e0"),
   384 => (x"87",x"e6",x"e9",x"4b"),
   385 => (x"c0",x"02",x"98",x"70"),
   386 => (x"48",x"c0",x"87",x"c5"),
   387 => (x"c2",x"87",x"f8",x"c3"),
   388 => (x"4c",x"bf",x"ce",x"ec"),
   389 => (x"5c",x"f7",x"f0",x"c2"),
   390 => (x"97",x"f3",x"e4",x"c2"),
   391 => (x"31",x"c8",x"49",x"bf"),
   392 => (x"97",x"f2",x"e4",x"c2"),
   393 => (x"49",x"a1",x"4a",x"bf"),
   394 => (x"97",x"f4",x"e4",x"c2"),
   395 => (x"32",x"d0",x"4a",x"bf"),
   396 => (x"c2",x"49",x"a1",x"72"),
   397 => (x"bf",x"97",x"f5",x"e4"),
   398 => (x"72",x"32",x"d8",x"4a"),
   399 => (x"66",x"c4",x"49",x"a1"),
   400 => (x"e3",x"f0",x"c2",x"91"),
   401 => (x"f0",x"c2",x"81",x"bf"),
   402 => (x"e4",x"c2",x"59",x"eb"),
   403 => (x"4a",x"bf",x"97",x"fb"),
   404 => (x"e4",x"c2",x"32",x"c8"),
   405 => (x"4b",x"bf",x"97",x"fa"),
   406 => (x"e4",x"c2",x"4a",x"a2"),
   407 => (x"4b",x"bf",x"97",x"fc"),
   408 => (x"a2",x"73",x"33",x"d0"),
   409 => (x"fd",x"e4",x"c2",x"4a"),
   410 => (x"cf",x"4b",x"bf",x"97"),
   411 => (x"73",x"33",x"d8",x"9b"),
   412 => (x"f0",x"c2",x"4a",x"a2"),
   413 => (x"f0",x"c2",x"5a",x"ef"),
   414 => (x"c2",x"4a",x"bf",x"eb"),
   415 => (x"c2",x"92",x"74",x"8a"),
   416 => (x"72",x"48",x"ef",x"f0"),
   417 => (x"ca",x"c1",x"78",x"a1"),
   418 => (x"e0",x"e4",x"c2",x"87"),
   419 => (x"c8",x"49",x"bf",x"97"),
   420 => (x"df",x"e4",x"c2",x"31"),
   421 => (x"a1",x"4a",x"bf",x"97"),
   422 => (x"de",x"ec",x"c2",x"49"),
   423 => (x"da",x"ec",x"c2",x"59"),
   424 => (x"31",x"c5",x"49",x"bf"),
   425 => (x"c9",x"81",x"ff",x"c7"),
   426 => (x"f7",x"f0",x"c2",x"29"),
   427 => (x"e5",x"e4",x"c2",x"59"),
   428 => (x"c8",x"4a",x"bf",x"97"),
   429 => (x"e4",x"e4",x"c2",x"32"),
   430 => (x"a2",x"4b",x"bf",x"97"),
   431 => (x"92",x"66",x"c4",x"4a"),
   432 => (x"f0",x"c2",x"82",x"6e"),
   433 => (x"f0",x"c2",x"5a",x"f3"),
   434 => (x"78",x"c0",x"48",x"eb"),
   435 => (x"48",x"e7",x"f0",x"c2"),
   436 => (x"c2",x"78",x"a1",x"72"),
   437 => (x"c2",x"48",x"f7",x"f0"),
   438 => (x"78",x"bf",x"eb",x"f0"),
   439 => (x"48",x"fb",x"f0",x"c2"),
   440 => (x"bf",x"ef",x"f0",x"c2"),
   441 => (x"d6",x"ec",x"c2",x"78"),
   442 => (x"c9",x"c0",x"02",x"bf"),
   443 => (x"c4",x"48",x"74",x"87"),
   444 => (x"c0",x"7e",x"70",x"30"),
   445 => (x"f0",x"c2",x"87",x"c9"),
   446 => (x"c4",x"48",x"bf",x"f3"),
   447 => (x"c2",x"7e",x"70",x"30"),
   448 => (x"6e",x"48",x"da",x"ec"),
   449 => (x"f8",x"48",x"c1",x"78"),
   450 => (x"26",x"4d",x"26",x"8e"),
   451 => (x"26",x"4b",x"26",x"4c"),
   452 => (x"5b",x"5e",x"0e",x"4f"),
   453 => (x"71",x"0e",x"5d",x"5c"),
   454 => (x"d6",x"ec",x"c2",x"4a"),
   455 => (x"87",x"cb",x"02",x"bf"),
   456 => (x"2b",x"c7",x"4b",x"72"),
   457 => (x"ff",x"c1",x"4c",x"72"),
   458 => (x"72",x"87",x"c9",x"9c"),
   459 => (x"72",x"2b",x"c8",x"4b"),
   460 => (x"9c",x"ff",x"c3",x"4c"),
   461 => (x"bf",x"e3",x"f0",x"c2"),
   462 => (x"c2",x"f5",x"c0",x"83"),
   463 => (x"d9",x"02",x"ab",x"bf"),
   464 => (x"c6",x"f5",x"c0",x"87"),
   465 => (x"ce",x"e4",x"c2",x"5b"),
   466 => (x"f0",x"49",x"73",x"1e"),
   467 => (x"86",x"c4",x"87",x"fd"),
   468 => (x"c5",x"05",x"98",x"70"),
   469 => (x"c0",x"48",x"c0",x"87"),
   470 => (x"ec",x"c2",x"87",x"e6"),
   471 => (x"d2",x"02",x"bf",x"d6"),
   472 => (x"c4",x"49",x"74",x"87"),
   473 => (x"ce",x"e4",x"c2",x"91"),
   474 => (x"cf",x"4d",x"69",x"81"),
   475 => (x"ff",x"ff",x"ff",x"ff"),
   476 => (x"74",x"87",x"cb",x"9d"),
   477 => (x"c2",x"91",x"c2",x"49"),
   478 => (x"9f",x"81",x"ce",x"e4"),
   479 => (x"48",x"75",x"4d",x"69"),
   480 => (x"0e",x"87",x"c6",x"fe"),
   481 => (x"5d",x"5c",x"5b",x"5e"),
   482 => (x"4d",x"71",x"1e",x"0e"),
   483 => (x"49",x"c1",x"1e",x"c0"),
   484 => (x"c4",x"87",x"d7",x"cf"),
   485 => (x"9c",x"4c",x"70",x"86"),
   486 => (x"87",x"c0",x"c1",x"02"),
   487 => (x"4a",x"de",x"ec",x"c2"),
   488 => (x"ea",x"e2",x"49",x"75"),
   489 => (x"02",x"98",x"70",x"87"),
   490 => (x"74",x"87",x"f1",x"c0"),
   491 => (x"cb",x"49",x"75",x"4a"),
   492 => (x"87",x"d0",x"e3",x"4b"),
   493 => (x"c0",x"02",x"98",x"70"),
   494 => (x"1e",x"c0",x"87",x"e2"),
   495 => (x"c7",x"02",x"9c",x"74"),
   496 => (x"48",x"a6",x"c4",x"87"),
   497 => (x"87",x"c5",x"78",x"c0"),
   498 => (x"c1",x"48",x"a6",x"c4"),
   499 => (x"49",x"66",x"c4",x"78"),
   500 => (x"c4",x"87",x"d7",x"ce"),
   501 => (x"9c",x"4c",x"70",x"86"),
   502 => (x"87",x"c0",x"ff",x"05"),
   503 => (x"fc",x"26",x"48",x"74"),
   504 => (x"5e",x"0e",x"87",x"e7"),
   505 => (x"0e",x"5d",x"5c",x"5b"),
   506 => (x"9b",x"4b",x"71",x"1e"),
   507 => (x"c0",x"87",x"c5",x"05"),
   508 => (x"87",x"e5",x"c1",x"48"),
   509 => (x"c0",x"4d",x"a3",x"c8"),
   510 => (x"02",x"66",x"d4",x"7d"),
   511 => (x"66",x"d4",x"87",x"c7"),
   512 => (x"c5",x"05",x"bf",x"97"),
   513 => (x"c1",x"48",x"c0",x"87"),
   514 => (x"66",x"d4",x"87",x"cf"),
   515 => (x"87",x"f3",x"fd",x"49"),
   516 => (x"02",x"9c",x"4c",x"70"),
   517 => (x"dc",x"87",x"c0",x"c1"),
   518 => (x"7d",x"69",x"49",x"a4"),
   519 => (x"c4",x"49",x"a4",x"da"),
   520 => (x"69",x"9f",x"4a",x"a3"),
   521 => (x"d6",x"ec",x"c2",x"7a"),
   522 => (x"87",x"d2",x"02",x"bf"),
   523 => (x"9f",x"49",x"a4",x"d4"),
   524 => (x"ff",x"c0",x"49",x"69"),
   525 => (x"48",x"71",x"99",x"ff"),
   526 => (x"7e",x"70",x"30",x"d0"),
   527 => (x"7e",x"c0",x"87",x"c2"),
   528 => (x"6a",x"48",x"49",x"6e"),
   529 => (x"c0",x"7a",x"70",x"80"),
   530 => (x"49",x"a3",x"cc",x"7b"),
   531 => (x"a3",x"d0",x"79",x"6a"),
   532 => (x"74",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"ec",x"fa",x"26",x"48"),
   535 => (x"5b",x"5e",x"0e",x"87"),
   536 => (x"71",x"0e",x"5d",x"5c"),
   537 => (x"c2",x"f5",x"c0",x"4c"),
   538 => (x"74",x"78",x"ff",x"48"),
   539 => (x"ca",x"c1",x"02",x"9c"),
   540 => (x"49",x"a4",x"c8",x"87"),
   541 => (x"c2",x"c1",x"02",x"69"),
   542 => (x"4a",x"66",x"d0",x"87"),
   543 => (x"d4",x"82",x"49",x"6c"),
   544 => (x"66",x"d0",x"5a",x"a6"),
   545 => (x"ec",x"c2",x"b9",x"4d"),
   546 => (x"ff",x"4a",x"bf",x"d2"),
   547 => (x"71",x"99",x"72",x"ba"),
   548 => (x"e4",x"c0",x"02",x"99"),
   549 => (x"4b",x"a4",x"c4",x"87"),
   550 => (x"f4",x"f9",x"49",x"6b"),
   551 => (x"c2",x"7b",x"70",x"87"),
   552 => (x"49",x"bf",x"ce",x"ec"),
   553 => (x"7c",x"71",x"81",x"6c"),
   554 => (x"ec",x"c2",x"b9",x"75"),
   555 => (x"ff",x"4a",x"bf",x"d2"),
   556 => (x"71",x"99",x"72",x"ba"),
   557 => (x"dc",x"ff",x"05",x"99"),
   558 => (x"f9",x"7c",x"75",x"87"),
   559 => (x"73",x"1e",x"87",x"cb"),
   560 => (x"9b",x"4b",x"71",x"1e"),
   561 => (x"c8",x"87",x"c7",x"02"),
   562 => (x"05",x"69",x"49",x"a3"),
   563 => (x"48",x"c0",x"87",x"c5"),
   564 => (x"c2",x"87",x"eb",x"c0"),
   565 => (x"4a",x"bf",x"e7",x"f0"),
   566 => (x"69",x"49",x"a3",x"c4"),
   567 => (x"c2",x"89",x"c2",x"49"),
   568 => (x"91",x"bf",x"ce",x"ec"),
   569 => (x"c2",x"4a",x"a2",x"71"),
   570 => (x"49",x"bf",x"d2",x"ec"),
   571 => (x"a2",x"71",x"99",x"6b"),
   572 => (x"1e",x"66",x"c8",x"4a"),
   573 => (x"d2",x"ea",x"49",x"72"),
   574 => (x"70",x"86",x"c4",x"87"),
   575 => (x"cc",x"f8",x"48",x"49"),
   576 => (x"5b",x"5e",x"0e",x"87"),
   577 => (x"1e",x"0e",x"5d",x"5c"),
   578 => (x"66",x"d4",x"4b",x"71"),
   579 => (x"73",x"2c",x"c9",x"4c"),
   580 => (x"cf",x"c1",x"02",x"9b"),
   581 => (x"49",x"a3",x"c8",x"87"),
   582 => (x"c7",x"c1",x"02",x"69"),
   583 => (x"4d",x"a3",x"d0",x"87"),
   584 => (x"c2",x"7d",x"66",x"d4"),
   585 => (x"49",x"bf",x"d2",x"ec"),
   586 => (x"4a",x"6b",x"b9",x"ff"),
   587 => (x"ac",x"71",x"7e",x"99"),
   588 => (x"c0",x"87",x"cd",x"03"),
   589 => (x"a3",x"cc",x"7d",x"7b"),
   590 => (x"49",x"a3",x"c4",x"4a"),
   591 => (x"87",x"c2",x"79",x"6a"),
   592 => (x"9c",x"74",x"8c",x"72"),
   593 => (x"49",x"87",x"dd",x"02"),
   594 => (x"fc",x"49",x"73",x"1e"),
   595 => (x"86",x"c4",x"87",x"cf"),
   596 => (x"c7",x"49",x"66",x"d4"),
   597 => (x"cb",x"02",x"99",x"ff"),
   598 => (x"ce",x"e4",x"c2",x"87"),
   599 => (x"fd",x"49",x"73",x"1e"),
   600 => (x"86",x"c4",x"87",x"dc"),
   601 => (x"87",x"e1",x"f6",x"26"),
   602 => (x"5c",x"5b",x"5e",x"0e"),
   603 => (x"86",x"f0",x"0e",x"5d"),
   604 => (x"c0",x"59",x"a6",x"d0"),
   605 => (x"cc",x"4b",x"66",x"e4"),
   606 => (x"87",x"ca",x"02",x"66"),
   607 => (x"70",x"80",x"c8",x"48"),
   608 => (x"05",x"bf",x"6e",x"7e"),
   609 => (x"48",x"c0",x"87",x"c5"),
   610 => (x"cc",x"87",x"ec",x"c3"),
   611 => (x"84",x"d0",x"4c",x"66"),
   612 => (x"a6",x"c4",x"49",x"73"),
   613 => (x"c4",x"78",x"6c",x"48"),
   614 => (x"80",x"c4",x"81",x"66"),
   615 => (x"c8",x"78",x"bf",x"6e"),
   616 => (x"c6",x"06",x"a9",x"66"),
   617 => (x"66",x"c4",x"49",x"87"),
   618 => (x"c0",x"4b",x"71",x"89"),
   619 => (x"c4",x"01",x"ab",x"b7"),
   620 => (x"c2",x"c3",x"48",x"87"),
   621 => (x"48",x"66",x"c4",x"87"),
   622 => (x"70",x"98",x"ff",x"c7"),
   623 => (x"c1",x"02",x"6e",x"7e"),
   624 => (x"c0",x"c8",x"87",x"c9"),
   625 => (x"71",x"89",x"6e",x"49"),
   626 => (x"ce",x"e4",x"c2",x"4a"),
   627 => (x"73",x"85",x"6e",x"4d"),
   628 => (x"c1",x"06",x"aa",x"b7"),
   629 => (x"49",x"72",x"4a",x"87"),
   630 => (x"80",x"66",x"c4",x"48"),
   631 => (x"8b",x"72",x"7c",x"70"),
   632 => (x"71",x"8a",x"c1",x"49"),
   633 => (x"87",x"d9",x"02",x"99"),
   634 => (x"48",x"66",x"e0",x"c0"),
   635 => (x"e0",x"c0",x"50",x"15"),
   636 => (x"80",x"c1",x"48",x"66"),
   637 => (x"58",x"a6",x"e4",x"c0"),
   638 => (x"8a",x"c1",x"49",x"72"),
   639 => (x"e7",x"05",x"99",x"71"),
   640 => (x"d0",x"1e",x"c1",x"87"),
   641 => (x"d4",x"f9",x"49",x"66"),
   642 => (x"c0",x"86",x"c4",x"87"),
   643 => (x"c1",x"06",x"ab",x"b7"),
   644 => (x"e0",x"c0",x"87",x"e3"),
   645 => (x"ff",x"c7",x"4d",x"66"),
   646 => (x"c0",x"06",x"ab",x"b7"),
   647 => (x"1e",x"75",x"87",x"e2"),
   648 => (x"fa",x"49",x"66",x"d0"),
   649 => (x"c0",x"c8",x"87",x"d8"),
   650 => (x"c8",x"48",x"6c",x"85"),
   651 => (x"7c",x"70",x"80",x"c0"),
   652 => (x"c1",x"8b",x"c0",x"c8"),
   653 => (x"49",x"66",x"d4",x"1e"),
   654 => (x"c8",x"87",x"e2",x"f8"),
   655 => (x"87",x"ee",x"c0",x"86"),
   656 => (x"1e",x"ce",x"e4",x"c2"),
   657 => (x"f9",x"49",x"66",x"d0"),
   658 => (x"86",x"c4",x"87",x"f4"),
   659 => (x"4a",x"ce",x"e4",x"c2"),
   660 => (x"6c",x"48",x"49",x"73"),
   661 => (x"73",x"7c",x"70",x"80"),
   662 => (x"71",x"8b",x"c1",x"49"),
   663 => (x"87",x"ce",x"02",x"99"),
   664 => (x"c1",x"7d",x"97",x"12"),
   665 => (x"c1",x"49",x"73",x"85"),
   666 => (x"05",x"99",x"71",x"8b"),
   667 => (x"b7",x"c0",x"87",x"f2"),
   668 => (x"e1",x"fe",x"01",x"ab"),
   669 => (x"f0",x"48",x"c1",x"87"),
   670 => (x"87",x"cd",x"f2",x"8e"),
   671 => (x"5c",x"5b",x"5e",x"0e"),
   672 => (x"4b",x"71",x"0e",x"5d"),
   673 => (x"87",x"c7",x"02",x"9b"),
   674 => (x"6d",x"4d",x"a3",x"c8"),
   675 => (x"ff",x"87",x"c5",x"05"),
   676 => (x"87",x"fd",x"c0",x"48"),
   677 => (x"6c",x"4c",x"a3",x"d0"),
   678 => (x"99",x"ff",x"c7",x"49"),
   679 => (x"6c",x"87",x"d8",x"05"),
   680 => (x"c1",x"87",x"c9",x"02"),
   681 => (x"f6",x"49",x"73",x"1e"),
   682 => (x"86",x"c4",x"87",x"f3"),
   683 => (x"1e",x"ce",x"e4",x"c2"),
   684 => (x"c9",x"f8",x"49",x"73"),
   685 => (x"6c",x"86",x"c4",x"87"),
   686 => (x"04",x"aa",x"6d",x"4a"),
   687 => (x"48",x"ff",x"87",x"c4"),
   688 => (x"a2",x"c1",x"87",x"cf"),
   689 => (x"c7",x"49",x"72",x"7c"),
   690 => (x"e4",x"c2",x"99",x"ff"),
   691 => (x"69",x"97",x"81",x"ce"),
   692 => (x"87",x"f5",x"f0",x"48"),
   693 => (x"71",x"1e",x"73",x"1e"),
   694 => (x"c0",x"02",x"9b",x"4b"),
   695 => (x"f0",x"c2",x"87",x"e4"),
   696 => (x"4a",x"73",x"5b",x"fb"),
   697 => (x"ec",x"c2",x"8a",x"c2"),
   698 => (x"92",x"49",x"bf",x"ce"),
   699 => (x"bf",x"e7",x"f0",x"c2"),
   700 => (x"c2",x"80",x"72",x"48"),
   701 => (x"71",x"58",x"ff",x"f0"),
   702 => (x"c2",x"30",x"c4",x"48"),
   703 => (x"c0",x"58",x"de",x"ec"),
   704 => (x"f0",x"c2",x"87",x"ed"),
   705 => (x"f0",x"c2",x"48",x"f7"),
   706 => (x"c2",x"78",x"bf",x"eb"),
   707 => (x"c2",x"48",x"fb",x"f0"),
   708 => (x"78",x"bf",x"ef",x"f0"),
   709 => (x"bf",x"d6",x"ec",x"c2"),
   710 => (x"c2",x"87",x"c9",x"02"),
   711 => (x"49",x"bf",x"ce",x"ec"),
   712 => (x"87",x"c7",x"31",x"c4"),
   713 => (x"bf",x"f3",x"f0",x"c2"),
   714 => (x"c2",x"31",x"c4",x"49"),
   715 => (x"ef",x"59",x"de",x"ec"),
   716 => (x"5e",x"0e",x"87",x"db"),
   717 => (x"71",x"0e",x"5c",x"5b"),
   718 => (x"72",x"4b",x"c0",x"4a"),
   719 => (x"e1",x"c0",x"02",x"9a"),
   720 => (x"49",x"a2",x"da",x"87"),
   721 => (x"c2",x"4b",x"69",x"9f"),
   722 => (x"02",x"bf",x"d6",x"ec"),
   723 => (x"a2",x"d4",x"87",x"cf"),
   724 => (x"49",x"69",x"9f",x"49"),
   725 => (x"ff",x"ff",x"c0",x"4c"),
   726 => (x"c2",x"34",x"d0",x"9c"),
   727 => (x"74",x"4c",x"c0",x"87"),
   728 => (x"49",x"73",x"b3",x"49"),
   729 => (x"ee",x"87",x"ed",x"fd"),
   730 => (x"5e",x"0e",x"87",x"e1"),
   731 => (x"0e",x"5d",x"5c",x"5b"),
   732 => (x"4a",x"71",x"86",x"f4"),
   733 => (x"9a",x"72",x"7e",x"c0"),
   734 => (x"c2",x"87",x"d8",x"02"),
   735 => (x"c0",x"48",x"ca",x"e4"),
   736 => (x"c2",x"e4",x"c2",x"78"),
   737 => (x"fb",x"f0",x"c2",x"48"),
   738 => (x"e4",x"c2",x"78",x"bf"),
   739 => (x"f0",x"c2",x"48",x"c6"),
   740 => (x"c2",x"78",x"bf",x"f7"),
   741 => (x"c0",x"48",x"eb",x"ec"),
   742 => (x"da",x"ec",x"c2",x"50"),
   743 => (x"e4",x"c2",x"49",x"bf"),
   744 => (x"71",x"4a",x"bf",x"ca"),
   745 => (x"c0",x"c4",x"03",x"aa"),
   746 => (x"cf",x"49",x"72",x"87"),
   747 => (x"e1",x"c0",x"05",x"99"),
   748 => (x"ce",x"e4",x"c2",x"87"),
   749 => (x"c2",x"e4",x"c2",x"1e"),
   750 => (x"e4",x"c2",x"49",x"bf"),
   751 => (x"a1",x"c1",x"48",x"c2"),
   752 => (x"df",x"ff",x"71",x"78"),
   753 => (x"86",x"c4",x"87",x"c5"),
   754 => (x"48",x"fe",x"f4",x"c0"),
   755 => (x"78",x"ce",x"e4",x"c2"),
   756 => (x"f4",x"c0",x"87",x"cc"),
   757 => (x"c0",x"48",x"bf",x"fe"),
   758 => (x"f5",x"c0",x"80",x"e0"),
   759 => (x"e4",x"c2",x"58",x"c2"),
   760 => (x"c1",x"48",x"bf",x"ca"),
   761 => (x"ce",x"e4",x"c2",x"80"),
   762 => (x"0d",x"3e",x"27",x"58"),
   763 => (x"97",x"bf",x"00",x"00"),
   764 => (x"02",x"9d",x"4d",x"bf"),
   765 => (x"c3",x"87",x"e2",x"c2"),
   766 => (x"c2",x"02",x"ad",x"e5"),
   767 => (x"f4",x"c0",x"87",x"db"),
   768 => (x"cb",x"4b",x"bf",x"fe"),
   769 => (x"4c",x"11",x"49",x"a3"),
   770 => (x"c1",x"05",x"ac",x"cf"),
   771 => (x"49",x"75",x"87",x"d2"),
   772 => (x"89",x"c1",x"99",x"df"),
   773 => (x"ec",x"c2",x"91",x"cd"),
   774 => (x"a3",x"c1",x"81",x"de"),
   775 => (x"c3",x"51",x"12",x"4a"),
   776 => (x"51",x"12",x"4a",x"a3"),
   777 => (x"12",x"4a",x"a3",x"c5"),
   778 => (x"4a",x"a3",x"c7",x"51"),
   779 => (x"a3",x"c9",x"51",x"12"),
   780 => (x"ce",x"51",x"12",x"4a"),
   781 => (x"51",x"12",x"4a",x"a3"),
   782 => (x"12",x"4a",x"a3",x"d0"),
   783 => (x"4a",x"a3",x"d2",x"51"),
   784 => (x"a3",x"d4",x"51",x"12"),
   785 => (x"d6",x"51",x"12",x"4a"),
   786 => (x"51",x"12",x"4a",x"a3"),
   787 => (x"12",x"4a",x"a3",x"d8"),
   788 => (x"4a",x"a3",x"dc",x"51"),
   789 => (x"a3",x"de",x"51",x"12"),
   790 => (x"c1",x"51",x"12",x"4a"),
   791 => (x"87",x"f9",x"c0",x"7e"),
   792 => (x"99",x"c8",x"49",x"74"),
   793 => (x"87",x"ea",x"c0",x"05"),
   794 => (x"99",x"d0",x"49",x"74"),
   795 => (x"dc",x"87",x"d0",x"05"),
   796 => (x"ca",x"c0",x"02",x"66"),
   797 => (x"dc",x"49",x"73",x"87"),
   798 => (x"98",x"70",x"0f",x"66"),
   799 => (x"6e",x"87",x"d3",x"02"),
   800 => (x"87",x"c6",x"c0",x"05"),
   801 => (x"48",x"de",x"ec",x"c2"),
   802 => (x"f4",x"c0",x"50",x"c0"),
   803 => (x"c2",x"48",x"bf",x"fe"),
   804 => (x"ec",x"c2",x"87",x"e7"),
   805 => (x"50",x"c0",x"48",x"eb"),
   806 => (x"da",x"ec",x"c2",x"7e"),
   807 => (x"e4",x"c2",x"49",x"bf"),
   808 => (x"71",x"4a",x"bf",x"ca"),
   809 => (x"c0",x"fc",x"04",x"aa"),
   810 => (x"fb",x"f0",x"c2",x"87"),
   811 => (x"c8",x"c0",x"05",x"bf"),
   812 => (x"d6",x"ec",x"c2",x"87"),
   813 => (x"fe",x"c1",x"02",x"bf"),
   814 => (x"c2",x"f5",x"c0",x"87"),
   815 => (x"c2",x"78",x"ff",x"48"),
   816 => (x"49",x"bf",x"c6",x"e4"),
   817 => (x"70",x"87",x"ca",x"e9"),
   818 => (x"ca",x"e4",x"c2",x"49"),
   819 => (x"48",x"a6",x"c4",x"59"),
   820 => (x"bf",x"c6",x"e4",x"c2"),
   821 => (x"d6",x"ec",x"c2",x"78"),
   822 => (x"d8",x"c0",x"02",x"bf"),
   823 => (x"49",x"66",x"c4",x"87"),
   824 => (x"ff",x"ff",x"ff",x"cf"),
   825 => (x"02",x"a9",x"99",x"f8"),
   826 => (x"c0",x"87",x"c5",x"c0"),
   827 => (x"87",x"e1",x"c0",x"4d"),
   828 => (x"dc",x"c0",x"4d",x"c1"),
   829 => (x"49",x"66",x"c4",x"87"),
   830 => (x"99",x"f8",x"ff",x"cf"),
   831 => (x"c8",x"c0",x"02",x"a9"),
   832 => (x"48",x"a6",x"c8",x"87"),
   833 => (x"c5",x"c0",x"78",x"c0"),
   834 => (x"48",x"a6",x"c8",x"87"),
   835 => (x"66",x"c8",x"78",x"c1"),
   836 => (x"05",x"9d",x"75",x"4d"),
   837 => (x"c4",x"87",x"e0",x"c0"),
   838 => (x"89",x"c2",x"49",x"66"),
   839 => (x"bf",x"ce",x"ec",x"c2"),
   840 => (x"f0",x"c2",x"91",x"4a"),
   841 => (x"c2",x"4a",x"bf",x"e7"),
   842 => (x"72",x"48",x"c2",x"e4"),
   843 => (x"e4",x"c2",x"78",x"a1"),
   844 => (x"78",x"c0",x"48",x"ca"),
   845 => (x"c0",x"87",x"e2",x"f9"),
   846 => (x"e7",x"8e",x"f4",x"48"),
   847 => (x"00",x"00",x"87",x"cb"),
   848 => (x"ff",x"ff",x"00",x"00"),
   849 => (x"0d",x"4e",x"ff",x"ff"),
   850 => (x"0d",x"57",x"00",x"00"),
   851 => (x"41",x"46",x"00",x"00"),
   852 => (x"20",x"32",x"33",x"54"),
   853 => (x"46",x"00",x"20",x"20"),
   854 => (x"36",x"31",x"54",x"41"),
   855 => (x"00",x"20",x"20",x"20"),
   856 => (x"c0",x"f1",x"c2",x"1e"),
   857 => (x"a8",x"dd",x"48",x"bf"),
   858 => (x"c0",x"87",x"c9",x"05"),
   859 => (x"70",x"87",x"ee",x"fe"),
   860 => (x"87",x"c8",x"4a",x"49"),
   861 => (x"c3",x"48",x"d4",x"ff"),
   862 => (x"4a",x"68",x"78",x"ff"),
   863 => (x"4f",x"26",x"48",x"72"),
   864 => (x"c0",x"f1",x"c2",x"1e"),
   865 => (x"a8",x"dd",x"48",x"bf"),
   866 => (x"c0",x"87",x"c6",x"05"),
   867 => (x"d9",x"87",x"fa",x"fd"),
   868 => (x"48",x"d4",x"ff",x"87"),
   869 => (x"ff",x"78",x"ff",x"c3"),
   870 => (x"e1",x"c8",x"48",x"d0"),
   871 => (x"48",x"d4",x"ff",x"78"),
   872 => (x"f0",x"c2",x"78",x"d4"),
   873 => (x"d4",x"ff",x"48",x"ff"),
   874 => (x"4f",x"26",x"50",x"bf"),
   875 => (x"48",x"d0",x"ff",x"1e"),
   876 => (x"26",x"78",x"e0",x"c0"),
   877 => (x"e7",x"fe",x"1e",x"4f"),
   878 => (x"99",x"49",x"70",x"87"),
   879 => (x"c0",x"87",x"c6",x"02"),
   880 => (x"f1",x"05",x"a9",x"fb"),
   881 => (x"26",x"48",x"71",x"87"),
   882 => (x"5b",x"5e",x"0e",x"4f"),
   883 => (x"4b",x"71",x"0e",x"5c"),
   884 => (x"cb",x"fe",x"4c",x"c0"),
   885 => (x"99",x"49",x"70",x"87"),
   886 => (x"87",x"f9",x"c0",x"02"),
   887 => (x"02",x"a9",x"ec",x"c0"),
   888 => (x"c0",x"87",x"f2",x"c0"),
   889 => (x"c0",x"02",x"a9",x"fb"),
   890 => (x"66",x"cc",x"87",x"eb"),
   891 => (x"c7",x"03",x"ac",x"b7"),
   892 => (x"02",x"66",x"d0",x"87"),
   893 => (x"53",x"71",x"87",x"c2"),
   894 => (x"c2",x"02",x"99",x"71"),
   895 => (x"fd",x"84",x"c1",x"87"),
   896 => (x"49",x"70",x"87",x"de"),
   897 => (x"87",x"cd",x"02",x"99"),
   898 => (x"02",x"a9",x"ec",x"c0"),
   899 => (x"fb",x"c0",x"87",x"c7"),
   900 => (x"d5",x"ff",x"05",x"a9"),
   901 => (x"02",x"66",x"d0",x"87"),
   902 => (x"97",x"c0",x"87",x"c3"),
   903 => (x"a9",x"ec",x"c0",x"7b"),
   904 => (x"74",x"87",x"c4",x"05"),
   905 => (x"74",x"87",x"c5",x"4a"),
   906 => (x"8a",x"0a",x"c0",x"4a"),
   907 => (x"87",x"c2",x"48",x"72"),
   908 => (x"4c",x"26",x"4d",x"26"),
   909 => (x"4f",x"26",x"4b",x"26"),
   910 => (x"87",x"e4",x"fc",x"1e"),
   911 => (x"f0",x"c0",x"49",x"70"),
   912 => (x"ca",x"04",x"a9",x"b7"),
   913 => (x"b7",x"f9",x"c0",x"87"),
   914 => (x"87",x"c3",x"01",x"a9"),
   915 => (x"c1",x"89",x"f0",x"c0"),
   916 => (x"04",x"a9",x"b7",x"c1"),
   917 => (x"da",x"c1",x"87",x"ca"),
   918 => (x"c3",x"01",x"a9",x"b7"),
   919 => (x"89",x"f7",x"c0",x"87"),
   920 => (x"4f",x"26",x"48",x"71"),
   921 => (x"5c",x"5b",x"5e",x"0e"),
   922 => (x"ff",x"4a",x"71",x"0e"),
   923 => (x"49",x"72",x"4c",x"d4"),
   924 => (x"70",x"87",x"ea",x"c0"),
   925 => (x"c2",x"02",x"9b",x"4b"),
   926 => (x"ff",x"8b",x"c1",x"87"),
   927 => (x"c5",x"c8",x"48",x"d0"),
   928 => (x"7c",x"d5",x"c1",x"78"),
   929 => (x"31",x"c6",x"49",x"73"),
   930 => (x"97",x"d2",x"e2",x"c2"),
   931 => (x"71",x"48",x"4a",x"bf"),
   932 => (x"ff",x"7c",x"70",x"b0"),
   933 => (x"78",x"c4",x"48",x"d0"),
   934 => (x"d5",x"fe",x"48",x"73"),
   935 => (x"5b",x"5e",x"0e",x"87"),
   936 => (x"f4",x"0e",x"5d",x"5c"),
   937 => (x"c4",x"4c",x"71",x"86"),
   938 => (x"78",x"c0",x"48",x"a6"),
   939 => (x"6e",x"7e",x"a4",x"c8"),
   940 => (x"c1",x"49",x"bf",x"97"),
   941 => (x"dd",x"05",x"a9",x"c1"),
   942 => (x"49",x"a4",x"c9",x"87"),
   943 => (x"c1",x"49",x"69",x"97"),
   944 => (x"d1",x"05",x"a9",x"d2"),
   945 => (x"49",x"a4",x"ca",x"87"),
   946 => (x"c1",x"49",x"69",x"97"),
   947 => (x"c5",x"05",x"a9",x"c3"),
   948 => (x"c2",x"48",x"df",x"87"),
   949 => (x"e7",x"fa",x"87",x"e1"),
   950 => (x"c0",x"4b",x"c0",x"87"),
   951 => (x"bf",x"97",x"fc",x"fd"),
   952 => (x"04",x"a9",x"c0",x"49"),
   953 => (x"cc",x"fb",x"87",x"cf"),
   954 => (x"c0",x"83",x"c1",x"87"),
   955 => (x"bf",x"97",x"fc",x"fd"),
   956 => (x"f1",x"06",x"ab",x"49"),
   957 => (x"fc",x"fd",x"c0",x"87"),
   958 => (x"cf",x"02",x"bf",x"97"),
   959 => (x"87",x"e0",x"f9",x"87"),
   960 => (x"02",x"99",x"49",x"70"),
   961 => (x"ec",x"c0",x"87",x"c6"),
   962 => (x"87",x"f1",x"05",x"a9"),
   963 => (x"cf",x"f9",x"4b",x"c0"),
   964 => (x"f9",x"4d",x"70",x"87"),
   965 => (x"a6",x"cc",x"87",x"ca"),
   966 => (x"87",x"c4",x"f9",x"58"),
   967 => (x"83",x"c1",x"4a",x"70"),
   968 => (x"49",x"bf",x"97",x"6e"),
   969 => (x"87",x"c7",x"02",x"ad"),
   970 => (x"05",x"ad",x"ff",x"c0"),
   971 => (x"c9",x"87",x"ea",x"c0"),
   972 => (x"69",x"97",x"49",x"a4"),
   973 => (x"a9",x"66",x"c8",x"49"),
   974 => (x"48",x"87",x"c7",x"02"),
   975 => (x"05",x"a8",x"ff",x"c0"),
   976 => (x"a4",x"ca",x"87",x"d7"),
   977 => (x"49",x"69",x"97",x"49"),
   978 => (x"87",x"c6",x"02",x"aa"),
   979 => (x"05",x"aa",x"ff",x"c0"),
   980 => (x"a6",x"c4",x"87",x"c7"),
   981 => (x"d3",x"78",x"c1",x"48"),
   982 => (x"ad",x"ec",x"c0",x"87"),
   983 => (x"c0",x"87",x"c6",x"02"),
   984 => (x"c7",x"05",x"ad",x"fb"),
   985 => (x"c4",x"4b",x"c0",x"87"),
   986 => (x"78",x"c1",x"48",x"a6"),
   987 => (x"fe",x"02",x"66",x"c4"),
   988 => (x"f7",x"f8",x"87",x"dc"),
   989 => (x"f4",x"48",x"73",x"87"),
   990 => (x"87",x"f4",x"fa",x"8e"),
   991 => (x"5b",x"5e",x"0e",x"00"),
   992 => (x"1e",x"0e",x"5d",x"5c"),
   993 => (x"4c",x"c0",x"4b",x"71"),
   994 => (x"c0",x"04",x"ab",x"4d"),
   995 => (x"fa",x"c0",x"87",x"e8"),
   996 => (x"9d",x"75",x"1e",x"dd"),
   997 => (x"c0",x"87",x"c4",x"02"),
   998 => (x"c1",x"87",x"c2",x"4a"),
   999 => (x"ef",x"49",x"72",x"4a"),
  1000 => (x"86",x"c4",x"87",x"c8"),
  1001 => (x"84",x"c1",x"7e",x"70"),
  1002 => (x"87",x"c2",x"05",x"6e"),
  1003 => (x"85",x"c1",x"4c",x"73"),
  1004 => (x"ff",x"06",x"ac",x"73"),
  1005 => (x"48",x"6e",x"87",x"d8"),
  1006 => (x"26",x"4d",x"26",x"26"),
  1007 => (x"26",x"4b",x"26",x"4c"),
  1008 => (x"5b",x"5e",x"0e",x"4f"),
  1009 => (x"1e",x"0e",x"5d",x"5c"),
  1010 => (x"de",x"49",x"4c",x"71"),
  1011 => (x"d9",x"f1",x"c2",x"91"),
  1012 => (x"97",x"85",x"71",x"4d"),
  1013 => (x"dd",x"c1",x"02",x"6d"),
  1014 => (x"c4",x"f1",x"c2",x"87"),
  1015 => (x"82",x"74",x"4a",x"bf"),
  1016 => (x"d8",x"fe",x"49",x"72"),
  1017 => (x"6e",x"7e",x"70",x"87"),
  1018 => (x"87",x"f3",x"c0",x"02"),
  1019 => (x"4b",x"cc",x"f1",x"c2"),
  1020 => (x"49",x"cb",x"4a",x"6e"),
  1021 => (x"87",x"f0",x"c2",x"ff"),
  1022 => (x"93",x"cb",x"4b",x"74"),
  1023 => (x"83",x"ee",x"e1",x"c1"),
  1024 => (x"c0",x"c1",x"83",x"c4"),
  1025 => (x"49",x"74",x"7b",x"fa"),
  1026 => (x"87",x"dc",x"cd",x"c1"),
  1027 => (x"f1",x"c2",x"7b",x"75"),
  1028 => (x"49",x"bf",x"97",x"d8"),
  1029 => (x"cc",x"f1",x"c2",x"1e"),
  1030 => (x"e6",x"e1",x"c1",x"49"),
  1031 => (x"74",x"86",x"c4",x"87"),
  1032 => (x"c3",x"cd",x"c1",x"49"),
  1033 => (x"c1",x"49",x"c0",x"87"),
  1034 => (x"c2",x"87",x"e2",x"ce"),
  1035 => (x"c0",x"48",x"c0",x"f1"),
  1036 => (x"dd",x"49",x"c1",x"78"),
  1037 => (x"fd",x"26",x"87",x"cf"),
  1038 => (x"6f",x"4c",x"87",x"ff"),
  1039 => (x"6e",x"69",x"64",x"61"),
  1040 => (x"2e",x"2e",x"2e",x"67"),
  1041 => (x"5b",x"5e",x"0e",x"00"),
  1042 => (x"4b",x"71",x"0e",x"5c"),
  1043 => (x"c4",x"f1",x"c2",x"4a"),
  1044 => (x"49",x"72",x"82",x"bf"),
  1045 => (x"70",x"87",x"e6",x"fc"),
  1046 => (x"c4",x"02",x"9c",x"4c"),
  1047 => (x"d1",x"eb",x"49",x"87"),
  1048 => (x"c4",x"f1",x"c2",x"87"),
  1049 => (x"c1",x"78",x"c0",x"48"),
  1050 => (x"87",x"d9",x"dc",x"49"),
  1051 => (x"0e",x"87",x"cc",x"fd"),
  1052 => (x"5d",x"5c",x"5b",x"5e"),
  1053 => (x"c2",x"86",x"f4",x"0e"),
  1054 => (x"c0",x"4d",x"ce",x"e4"),
  1055 => (x"48",x"a6",x"c4",x"4c"),
  1056 => (x"f1",x"c2",x"78",x"c0"),
  1057 => (x"c0",x"49",x"bf",x"c4"),
  1058 => (x"c1",x"c1",x"06",x"a9"),
  1059 => (x"ce",x"e4",x"c2",x"87"),
  1060 => (x"c0",x"02",x"98",x"48"),
  1061 => (x"fa",x"c0",x"87",x"f8"),
  1062 => (x"66",x"c8",x"1e",x"dd"),
  1063 => (x"c4",x"87",x"c7",x"02"),
  1064 => (x"78",x"c0",x"48",x"a6"),
  1065 => (x"a6",x"c4",x"87",x"c5"),
  1066 => (x"c4",x"78",x"c1",x"48"),
  1067 => (x"f9",x"ea",x"49",x"66"),
  1068 => (x"70",x"86",x"c4",x"87"),
  1069 => (x"c4",x"84",x"c1",x"4d"),
  1070 => (x"80",x"c1",x"48",x"66"),
  1071 => (x"c2",x"58",x"a6",x"c8"),
  1072 => (x"49",x"bf",x"c4",x"f1"),
  1073 => (x"87",x"c6",x"03",x"ac"),
  1074 => (x"ff",x"05",x"9d",x"75"),
  1075 => (x"4c",x"c0",x"87",x"c8"),
  1076 => (x"c3",x"02",x"9d",x"75"),
  1077 => (x"fa",x"c0",x"87",x"e0"),
  1078 => (x"66",x"c8",x"1e",x"dd"),
  1079 => (x"cc",x"87",x"c7",x"02"),
  1080 => (x"78",x"c0",x"48",x"a6"),
  1081 => (x"a6",x"cc",x"87",x"c5"),
  1082 => (x"cc",x"78",x"c1",x"48"),
  1083 => (x"f9",x"e9",x"49",x"66"),
  1084 => (x"70",x"86",x"c4",x"87"),
  1085 => (x"c2",x"02",x"6e",x"7e"),
  1086 => (x"49",x"6e",x"87",x"e9"),
  1087 => (x"69",x"97",x"81",x"cb"),
  1088 => (x"02",x"99",x"d0",x"49"),
  1089 => (x"c1",x"87",x"d6",x"c1"),
  1090 => (x"74",x"4a",x"c5",x"c1"),
  1091 => (x"c1",x"91",x"cb",x"49"),
  1092 => (x"72",x"81",x"ee",x"e1"),
  1093 => (x"c3",x"81",x"c8",x"79"),
  1094 => (x"49",x"74",x"51",x"ff"),
  1095 => (x"f1",x"c2",x"91",x"de"),
  1096 => (x"85",x"71",x"4d",x"d9"),
  1097 => (x"7d",x"97",x"c1",x"c2"),
  1098 => (x"c0",x"49",x"a5",x"c1"),
  1099 => (x"ec",x"c2",x"51",x"e0"),
  1100 => (x"02",x"bf",x"97",x"de"),
  1101 => (x"84",x"c1",x"87",x"d2"),
  1102 => (x"c2",x"4b",x"a5",x"c2"),
  1103 => (x"db",x"4a",x"de",x"ec"),
  1104 => (x"e3",x"fd",x"fe",x"49"),
  1105 => (x"87",x"db",x"c1",x"87"),
  1106 => (x"c0",x"49",x"a5",x"cd"),
  1107 => (x"c2",x"84",x"c1",x"51"),
  1108 => (x"4a",x"6e",x"4b",x"a5"),
  1109 => (x"fd",x"fe",x"49",x"cb"),
  1110 => (x"c6",x"c1",x"87",x"ce"),
  1111 => (x"c1",x"ff",x"c0",x"87"),
  1112 => (x"cb",x"49",x"74",x"4a"),
  1113 => (x"ee",x"e1",x"c1",x"91"),
  1114 => (x"c2",x"79",x"72",x"81"),
  1115 => (x"bf",x"97",x"de",x"ec"),
  1116 => (x"74",x"87",x"d8",x"02"),
  1117 => (x"c1",x"91",x"de",x"49"),
  1118 => (x"d9",x"f1",x"c2",x"84"),
  1119 => (x"c2",x"83",x"71",x"4b"),
  1120 => (x"dd",x"4a",x"de",x"ec"),
  1121 => (x"df",x"fc",x"fe",x"49"),
  1122 => (x"74",x"87",x"d8",x"87"),
  1123 => (x"c2",x"93",x"de",x"4b"),
  1124 => (x"cb",x"83",x"d9",x"f1"),
  1125 => (x"51",x"c0",x"49",x"a3"),
  1126 => (x"6e",x"73",x"84",x"c1"),
  1127 => (x"fe",x"49",x"cb",x"4a"),
  1128 => (x"c4",x"87",x"c5",x"fc"),
  1129 => (x"80",x"c1",x"48",x"66"),
  1130 => (x"c7",x"58",x"a6",x"c8"),
  1131 => (x"c5",x"c0",x"03",x"ac"),
  1132 => (x"fc",x"05",x"6e",x"87"),
  1133 => (x"48",x"74",x"87",x"e0"),
  1134 => (x"fc",x"f7",x"8e",x"f4"),
  1135 => (x"1e",x"73",x"1e",x"87"),
  1136 => (x"cb",x"49",x"4b",x"71"),
  1137 => (x"ee",x"e1",x"c1",x"91"),
  1138 => (x"4a",x"a1",x"c8",x"81"),
  1139 => (x"48",x"d2",x"e2",x"c2"),
  1140 => (x"a1",x"c9",x"50",x"12"),
  1141 => (x"fc",x"fd",x"c0",x"4a"),
  1142 => (x"ca",x"50",x"12",x"48"),
  1143 => (x"d8",x"f1",x"c2",x"81"),
  1144 => (x"c2",x"50",x"11",x"48"),
  1145 => (x"bf",x"97",x"d8",x"f1"),
  1146 => (x"49",x"c0",x"1e",x"49"),
  1147 => (x"87",x"d3",x"da",x"c1"),
  1148 => (x"48",x"c0",x"f1",x"c2"),
  1149 => (x"49",x"c1",x"78",x"de"),
  1150 => (x"26",x"87",x"ca",x"d6"),
  1151 => (x"1e",x"87",x"fe",x"f6"),
  1152 => (x"cb",x"49",x"4a",x"71"),
  1153 => (x"ee",x"e1",x"c1",x"91"),
  1154 => (x"11",x"81",x"c8",x"81"),
  1155 => (x"c4",x"f1",x"c2",x"48"),
  1156 => (x"c4",x"f1",x"c2",x"58"),
  1157 => (x"c1",x"78",x"c0",x"48"),
  1158 => (x"87",x"e9",x"d5",x"49"),
  1159 => (x"c0",x"1e",x"4f",x"26"),
  1160 => (x"e8",x"c6",x"c1",x"49"),
  1161 => (x"1e",x"4f",x"26",x"87"),
  1162 => (x"d2",x"02",x"99",x"71"),
  1163 => (x"c3",x"e3",x"c1",x"87"),
  1164 => (x"f7",x"50",x"c0",x"48"),
  1165 => (x"ff",x"c7",x"c1",x"80"),
  1166 => (x"e7",x"e1",x"c1",x"40"),
  1167 => (x"c1",x"87",x"ce",x"78"),
  1168 => (x"c1",x"48",x"ff",x"e2"),
  1169 => (x"fc",x"78",x"e0",x"e1"),
  1170 => (x"de",x"c8",x"c1",x"80"),
  1171 => (x"0e",x"4f",x"26",x"78"),
  1172 => (x"0e",x"5c",x"5b",x"5e"),
  1173 => (x"cb",x"4a",x"4c",x"71"),
  1174 => (x"ee",x"e1",x"c1",x"92"),
  1175 => (x"49",x"a2",x"c8",x"82"),
  1176 => (x"97",x"4b",x"a2",x"c9"),
  1177 => (x"97",x"1e",x"4b",x"6b"),
  1178 => (x"ca",x"1e",x"49",x"69"),
  1179 => (x"c0",x"49",x"12",x"82"),
  1180 => (x"c0",x"87",x"c9",x"e7"),
  1181 => (x"87",x"cd",x"d4",x"49"),
  1182 => (x"c3",x"c1",x"49",x"74"),
  1183 => (x"8e",x"f8",x"87",x"ea"),
  1184 => (x"1e",x"87",x"f8",x"f4"),
  1185 => (x"4b",x"71",x"1e",x"73"),
  1186 => (x"87",x"c3",x"ff",x"49"),
  1187 => (x"fe",x"fe",x"49",x"73"),
  1188 => (x"87",x"e9",x"f4",x"87"),
  1189 => (x"71",x"1e",x"73",x"1e"),
  1190 => (x"4a",x"a3",x"c6",x"4b"),
  1191 => (x"c1",x"87",x"db",x"02"),
  1192 => (x"87",x"d6",x"02",x"8a"),
  1193 => (x"da",x"c1",x"02",x"8a"),
  1194 => (x"c0",x"02",x"8a",x"87"),
  1195 => (x"02",x"8a",x"87",x"fc"),
  1196 => (x"8a",x"87",x"e1",x"c0"),
  1197 => (x"c1",x"87",x"cb",x"02"),
  1198 => (x"49",x"c7",x"87",x"db"),
  1199 => (x"c1",x"87",x"c0",x"fd"),
  1200 => (x"f1",x"c2",x"87",x"de"),
  1201 => (x"c1",x"02",x"bf",x"c4"),
  1202 => (x"c1",x"48",x"87",x"cb"),
  1203 => (x"c8",x"f1",x"c2",x"88"),
  1204 => (x"87",x"c1",x"c1",x"58"),
  1205 => (x"bf",x"c8",x"f1",x"c2"),
  1206 => (x"87",x"f9",x"c0",x"02"),
  1207 => (x"bf",x"c4",x"f1",x"c2"),
  1208 => (x"c2",x"80",x"c1",x"48"),
  1209 => (x"c0",x"58",x"c8",x"f1"),
  1210 => (x"f1",x"c2",x"87",x"eb"),
  1211 => (x"c6",x"49",x"bf",x"c4"),
  1212 => (x"c8",x"f1",x"c2",x"89"),
  1213 => (x"a9",x"b7",x"c0",x"59"),
  1214 => (x"c2",x"87",x"da",x"03"),
  1215 => (x"c0",x"48",x"c4",x"f1"),
  1216 => (x"c2",x"87",x"d2",x"78"),
  1217 => (x"02",x"bf",x"c8",x"f1"),
  1218 => (x"f1",x"c2",x"87",x"cb"),
  1219 => (x"c6",x"48",x"bf",x"c4"),
  1220 => (x"c8",x"f1",x"c2",x"80"),
  1221 => (x"d1",x"49",x"c0",x"58"),
  1222 => (x"49",x"73",x"87",x"eb"),
  1223 => (x"87",x"c8",x"c1",x"c1"),
  1224 => (x"1e",x"87",x"da",x"f2"),
  1225 => (x"4b",x"71",x"1e",x"73"),
  1226 => (x"48",x"c0",x"f1",x"c2"),
  1227 => (x"49",x"c0",x"78",x"dd"),
  1228 => (x"73",x"87",x"d2",x"d1"),
  1229 => (x"ef",x"c0",x"c1",x"49"),
  1230 => (x"87",x"c1",x"f2",x"87"),
  1231 => (x"5c",x"5b",x"5e",x"0e"),
  1232 => (x"cc",x"4c",x"71",x"0e"),
  1233 => (x"4b",x"74",x"1e",x"66"),
  1234 => (x"e1",x"c1",x"93",x"cb"),
  1235 => (x"a3",x"c4",x"83",x"ee"),
  1236 => (x"fe",x"49",x"6a",x"4a"),
  1237 => (x"c1",x"87",x"e1",x"f5"),
  1238 => (x"c8",x"7b",x"fd",x"c6"),
  1239 => (x"66",x"d4",x"49",x"a3"),
  1240 => (x"49",x"a3",x"c9",x"51"),
  1241 => (x"ca",x"51",x"66",x"d8"),
  1242 => (x"66",x"dc",x"49",x"a3"),
  1243 => (x"ca",x"f1",x"26",x"51"),
  1244 => (x"5b",x"5e",x"0e",x"87"),
  1245 => (x"ff",x"0e",x"5d",x"5c"),
  1246 => (x"a6",x"dc",x"86",x"cc"),
  1247 => (x"48",x"a6",x"c8",x"59"),
  1248 => (x"80",x"c4",x"78",x"c0"),
  1249 => (x"78",x"66",x"c8",x"c1"),
  1250 => (x"78",x"c1",x"80",x"c4"),
  1251 => (x"78",x"c1",x"80",x"c4"),
  1252 => (x"48",x"c8",x"f1",x"c2"),
  1253 => (x"f1",x"c2",x"78",x"c1"),
  1254 => (x"de",x"48",x"bf",x"c0"),
  1255 => (x"87",x"cb",x"05",x"a8"),
  1256 => (x"70",x"87",x"cc",x"f3"),
  1257 => (x"59",x"a6",x"cc",x"49"),
  1258 => (x"e7",x"87",x"d6",x"ce"),
  1259 => (x"c4",x"e8",x"87",x"d2"),
  1260 => (x"87",x"ec",x"e6",x"87"),
  1261 => (x"fb",x"c0",x"4c",x"70"),
  1262 => (x"d8",x"c1",x"02",x"ac"),
  1263 => (x"05",x"66",x"d8",x"87"),
  1264 => (x"c0",x"87",x"ca",x"c1"),
  1265 => (x"1e",x"c1",x"1e",x"1e"),
  1266 => (x"1e",x"e1",x"e3",x"c1"),
  1267 => (x"eb",x"fd",x"49",x"c0"),
  1268 => (x"c0",x"86",x"d0",x"87"),
  1269 => (x"d9",x"02",x"ac",x"fb"),
  1270 => (x"66",x"c4",x"c1",x"87"),
  1271 => (x"6a",x"82",x"c4",x"4a"),
  1272 => (x"74",x"81",x"c7",x"49"),
  1273 => (x"d8",x"1e",x"c1",x"51"),
  1274 => (x"c8",x"49",x"6a",x"1e"),
  1275 => (x"87",x"d9",x"e7",x"81"),
  1276 => (x"c8",x"c1",x"86",x"c8"),
  1277 => (x"a8",x"c0",x"48",x"66"),
  1278 => (x"c8",x"87",x"c7",x"01"),
  1279 => (x"78",x"c1",x"48",x"a6"),
  1280 => (x"c8",x"c1",x"87",x"ce"),
  1281 => (x"88",x"c1",x"48",x"66"),
  1282 => (x"c3",x"58",x"a6",x"d0"),
  1283 => (x"87",x"e5",x"e6",x"87"),
  1284 => (x"c2",x"48",x"a6",x"d0"),
  1285 => (x"02",x"9c",x"74",x"78"),
  1286 => (x"c8",x"87",x"e2",x"cc"),
  1287 => (x"cc",x"c1",x"48",x"66"),
  1288 => (x"cc",x"03",x"a8",x"66"),
  1289 => (x"a6",x"dc",x"87",x"d7"),
  1290 => (x"e4",x"78",x"c0",x"48"),
  1291 => (x"4c",x"70",x"87",x"f2"),
  1292 => (x"dd",x"48",x"66",x"d8"),
  1293 => (x"87",x"c6",x"05",x"a8"),
  1294 => (x"d8",x"48",x"a6",x"dc"),
  1295 => (x"d0",x"c1",x"78",x"66"),
  1296 => (x"e8",x"c0",x"05",x"ac"),
  1297 => (x"87",x"d8",x"e4",x"87"),
  1298 => (x"70",x"87",x"d5",x"e4"),
  1299 => (x"ac",x"ec",x"c0",x"4c"),
  1300 => (x"e5",x"87",x"c5",x"05"),
  1301 => (x"4c",x"70",x"87",x"df"),
  1302 => (x"05",x"ac",x"d0",x"c1"),
  1303 => (x"66",x"d4",x"87",x"c8"),
  1304 => (x"d8",x"80",x"c1",x"48"),
  1305 => (x"d0",x"c1",x"58",x"a6"),
  1306 => (x"d8",x"ff",x"02",x"ac"),
  1307 => (x"a6",x"e0",x"c0",x"87"),
  1308 => (x"78",x"66",x"d8",x"48"),
  1309 => (x"c0",x"48",x"66",x"dc"),
  1310 => (x"05",x"a8",x"66",x"e0"),
  1311 => (x"c4",x"87",x"d0",x"ca"),
  1312 => (x"f0",x"c0",x"48",x"a6"),
  1313 => (x"80",x"e0",x"c0",x"78"),
  1314 => (x"c4",x"78",x"66",x"d0"),
  1315 => (x"c4",x"78",x"c0",x"80"),
  1316 => (x"74",x"78",x"c0",x"80"),
  1317 => (x"8d",x"fb",x"c0",x"4d"),
  1318 => (x"87",x"cc",x"c9",x"02"),
  1319 => (x"db",x"02",x"8d",x"c9"),
  1320 => (x"02",x"8d",x"c2",x"87"),
  1321 => (x"c9",x"87",x"cd",x"c1"),
  1322 => (x"d1",x"c4",x"02",x"8d"),
  1323 => (x"02",x"8d",x"c4",x"87"),
  1324 => (x"c1",x"87",x"ce",x"c1"),
  1325 => (x"c5",x"c4",x"02",x"8d"),
  1326 => (x"87",x"e6",x"c8",x"87"),
  1327 => (x"cb",x"49",x"66",x"c8"),
  1328 => (x"66",x"c4",x"c1",x"91"),
  1329 => (x"4a",x"a1",x"c4",x"81"),
  1330 => (x"1e",x"71",x"7e",x"6a"),
  1331 => (x"48",x"f8",x"dd",x"c1"),
  1332 => (x"cc",x"49",x"66",x"c4"),
  1333 => (x"41",x"20",x"4a",x"a1"),
  1334 => (x"ff",x"05",x"aa",x"71"),
  1335 => (x"51",x"10",x"87",x"f8"),
  1336 => (x"cc",x"c1",x"49",x"26"),
  1337 => (x"cc",x"e3",x"79",x"e3"),
  1338 => (x"c0",x"4c",x"70",x"87"),
  1339 => (x"c1",x"48",x"a6",x"ec"),
  1340 => (x"87",x"f4",x"c7",x"78"),
  1341 => (x"c0",x"48",x"a6",x"c4"),
  1342 => (x"48",x"66",x"d0",x"78"),
  1343 => (x"a6",x"d4",x"80",x"c1"),
  1344 => (x"87",x"dc",x"e1",x"58"),
  1345 => (x"ec",x"c0",x"4c",x"70"),
  1346 => (x"87",x"d4",x"02",x"ac"),
  1347 => (x"c0",x"02",x"66",x"c4"),
  1348 => (x"a6",x"c8",x"87",x"c5"),
  1349 => (x"74",x"87",x"c9",x"5c"),
  1350 => (x"88",x"f0",x"c0",x"48"),
  1351 => (x"58",x"a6",x"e8",x"c0"),
  1352 => (x"02",x"ac",x"ec",x"c0"),
  1353 => (x"f7",x"e0",x"87",x"cc"),
  1354 => (x"c0",x"4c",x"70",x"87"),
  1355 => (x"ff",x"05",x"ac",x"ec"),
  1356 => (x"66",x"c4",x"87",x"f4"),
  1357 => (x"49",x"66",x"d8",x"1e"),
  1358 => (x"66",x"ec",x"c0",x"1e"),
  1359 => (x"e1",x"e3",x"c1",x"1e"),
  1360 => (x"49",x"66",x"d8",x"1e"),
  1361 => (x"c0",x"87",x"f5",x"f7"),
  1362 => (x"c0",x"1e",x"ca",x"1e"),
  1363 => (x"cb",x"49",x"66",x"e0"),
  1364 => (x"66",x"dc",x"c1",x"91"),
  1365 => (x"48",x"a6",x"d8",x"81"),
  1366 => (x"d8",x"78",x"a1",x"c4"),
  1367 => (x"e1",x"49",x"bf",x"66"),
  1368 => (x"86",x"d8",x"87",x"e7"),
  1369 => (x"06",x"a8",x"b7",x"c0"),
  1370 => (x"c1",x"87",x"ca",x"c1"),
  1371 => (x"c8",x"1e",x"de",x"1e"),
  1372 => (x"e1",x"49",x"bf",x"66"),
  1373 => (x"86",x"c8",x"87",x"d3"),
  1374 => (x"c0",x"48",x"49",x"70"),
  1375 => (x"e8",x"c0",x"88",x"08"),
  1376 => (x"b7",x"c0",x"58",x"a6"),
  1377 => (x"ec",x"c0",x"06",x"a8"),
  1378 => (x"66",x"e4",x"c0",x"87"),
  1379 => (x"a8",x"b7",x"dd",x"48"),
  1380 => (x"87",x"e1",x"c0",x"03"),
  1381 => (x"c0",x"49",x"bf",x"6e"),
  1382 => (x"c0",x"81",x"66",x"e4"),
  1383 => (x"e4",x"c0",x"51",x"e0"),
  1384 => (x"81",x"c1",x"49",x"66"),
  1385 => (x"c2",x"81",x"bf",x"6e"),
  1386 => (x"e4",x"c0",x"51",x"c1"),
  1387 => (x"81",x"c2",x"49",x"66"),
  1388 => (x"c0",x"81",x"bf",x"6e"),
  1389 => (x"a6",x"ec",x"c0",x"51"),
  1390 => (x"c4",x"78",x"c1",x"48"),
  1391 => (x"f7",x"e1",x"87",x"ea"),
  1392 => (x"a6",x"e8",x"c0",x"87"),
  1393 => (x"87",x"f0",x"e1",x"58"),
  1394 => (x"58",x"a6",x"f0",x"c0"),
  1395 => (x"05",x"a8",x"ec",x"c0"),
  1396 => (x"a6",x"87",x"c9",x"c0"),
  1397 => (x"66",x"e4",x"c0",x"48"),
  1398 => (x"87",x"c4",x"c0",x"78"),
  1399 => (x"87",x"c0",x"de",x"ff"),
  1400 => (x"cb",x"49",x"66",x"c8"),
  1401 => (x"66",x"c4",x"c1",x"91"),
  1402 => (x"c8",x"80",x"71",x"48"),
  1403 => (x"66",x"c4",x"58",x"a6"),
  1404 => (x"c4",x"82",x"c8",x"4a"),
  1405 => (x"81",x"ca",x"49",x"66"),
  1406 => (x"51",x"66",x"e4",x"c0"),
  1407 => (x"49",x"66",x"ec",x"c0"),
  1408 => (x"e4",x"c0",x"81",x"c1"),
  1409 => (x"48",x"c1",x"89",x"66"),
  1410 => (x"49",x"70",x"30",x"71"),
  1411 => (x"97",x"71",x"89",x"c1"),
  1412 => (x"f5",x"f4",x"c2",x"7a"),
  1413 => (x"e4",x"c0",x"49",x"bf"),
  1414 => (x"6a",x"97",x"29",x"66"),
  1415 => (x"98",x"71",x"48",x"4a"),
  1416 => (x"58",x"a6",x"f4",x"c0"),
  1417 => (x"c4",x"49",x"66",x"c4"),
  1418 => (x"c0",x"7e",x"69",x"81"),
  1419 => (x"dc",x"48",x"66",x"e0"),
  1420 => (x"c0",x"02",x"a8",x"66"),
  1421 => (x"a6",x"dc",x"87",x"c8"),
  1422 => (x"c0",x"78",x"c0",x"48"),
  1423 => (x"a6",x"dc",x"87",x"c5"),
  1424 => (x"dc",x"78",x"c1",x"48"),
  1425 => (x"e0",x"c0",x"1e",x"66"),
  1426 => (x"49",x"66",x"c8",x"1e"),
  1427 => (x"87",x"f9",x"dd",x"ff"),
  1428 => (x"4c",x"70",x"86",x"c8"),
  1429 => (x"06",x"ac",x"b7",x"c0"),
  1430 => (x"6e",x"87",x"d6",x"c1"),
  1431 => (x"70",x"80",x"74",x"48"),
  1432 => (x"49",x"e0",x"c0",x"7e"),
  1433 => (x"4b",x"6e",x"89",x"74"),
  1434 => (x"4a",x"f5",x"dd",x"c1"),
  1435 => (x"f7",x"e8",x"fe",x"71"),
  1436 => (x"c2",x"48",x"6e",x"87"),
  1437 => (x"c0",x"7e",x"70",x"80"),
  1438 => (x"c1",x"48",x"66",x"e8"),
  1439 => (x"a6",x"ec",x"c0",x"80"),
  1440 => (x"66",x"f0",x"c0",x"58"),
  1441 => (x"70",x"81",x"c1",x"49"),
  1442 => (x"c5",x"c0",x"02",x"a9"),
  1443 => (x"c0",x"4d",x"c0",x"87"),
  1444 => (x"4d",x"c1",x"87",x"c2"),
  1445 => (x"a4",x"c2",x"1e",x"75"),
  1446 => (x"48",x"e0",x"c0",x"49"),
  1447 => (x"49",x"70",x"88",x"71"),
  1448 => (x"49",x"66",x"c8",x"1e"),
  1449 => (x"87",x"e1",x"dc",x"ff"),
  1450 => (x"b7",x"c0",x"86",x"c8"),
  1451 => (x"c6",x"ff",x"01",x"a8"),
  1452 => (x"66",x"e8",x"c0",x"87"),
  1453 => (x"87",x"d3",x"c0",x"02"),
  1454 => (x"c9",x"49",x"66",x"c4"),
  1455 => (x"66",x"e8",x"c0",x"81"),
  1456 => (x"48",x"66",x"c4",x"51"),
  1457 => (x"78",x"cf",x"c9",x"c1"),
  1458 => (x"c4",x"87",x"ce",x"c0"),
  1459 => (x"81",x"c9",x"49",x"66"),
  1460 => (x"66",x"c4",x"51",x"c2"),
  1461 => (x"c3",x"ca",x"c1",x"48"),
  1462 => (x"a6",x"ec",x"c0",x"78"),
  1463 => (x"c0",x"78",x"c1",x"48"),
  1464 => (x"db",x"ff",x"87",x"c6"),
  1465 => (x"4c",x"70",x"87",x"cf"),
  1466 => (x"02",x"66",x"ec",x"c0"),
  1467 => (x"c8",x"87",x"f5",x"c0"),
  1468 => (x"66",x"cc",x"48",x"66"),
  1469 => (x"cb",x"c0",x"04",x"a8"),
  1470 => (x"48",x"66",x"c8",x"87"),
  1471 => (x"a6",x"cc",x"80",x"c1"),
  1472 => (x"87",x"e0",x"c0",x"58"),
  1473 => (x"c1",x"48",x"66",x"cc"),
  1474 => (x"58",x"a6",x"d0",x"88"),
  1475 => (x"c1",x"87",x"d5",x"c0"),
  1476 => (x"c0",x"05",x"ac",x"c6"),
  1477 => (x"66",x"d0",x"87",x"c8"),
  1478 => (x"d4",x"80",x"c1",x"48"),
  1479 => (x"da",x"ff",x"58",x"a6"),
  1480 => (x"4c",x"70",x"87",x"d3"),
  1481 => (x"c1",x"48",x"66",x"d4"),
  1482 => (x"58",x"a6",x"d8",x"80"),
  1483 => (x"c0",x"02",x"9c",x"74"),
  1484 => (x"66",x"c8",x"87",x"cb"),
  1485 => (x"66",x"cc",x"c1",x"48"),
  1486 => (x"e9",x"f3",x"04",x"a8"),
  1487 => (x"eb",x"d9",x"ff",x"87"),
  1488 => (x"48",x"66",x"c8",x"87"),
  1489 => (x"c0",x"03",x"a8",x"c7"),
  1490 => (x"f1",x"c2",x"87",x"e5"),
  1491 => (x"78",x"c0",x"48",x"c8"),
  1492 => (x"cb",x"49",x"66",x"c8"),
  1493 => (x"66",x"c4",x"c1",x"91"),
  1494 => (x"4a",x"a1",x"c4",x"81"),
  1495 => (x"52",x"c0",x"4a",x"6a"),
  1496 => (x"48",x"66",x"c8",x"79"),
  1497 => (x"a6",x"cc",x"80",x"c1"),
  1498 => (x"04",x"a8",x"c7",x"58"),
  1499 => (x"ff",x"87",x"db",x"ff"),
  1500 => (x"c4",x"e1",x"8e",x"cc"),
  1501 => (x"00",x"20",x"3a",x"87"),
  1502 => (x"20",x"50",x"49",x"44"),
  1503 => (x"74",x"69",x"77",x"53"),
  1504 => (x"73",x"65",x"68",x"63"),
  1505 => (x"1e",x"73",x"1e",x"00"),
  1506 => (x"02",x"9b",x"4b",x"71"),
  1507 => (x"f1",x"c2",x"87",x"c6"),
  1508 => (x"78",x"c0",x"48",x"c4"),
  1509 => (x"f1",x"c2",x"1e",x"c7"),
  1510 => (x"1e",x"49",x"bf",x"c4"),
  1511 => (x"1e",x"ee",x"e1",x"c1"),
  1512 => (x"bf",x"c0",x"f1",x"c2"),
  1513 => (x"87",x"c9",x"ef",x"49"),
  1514 => (x"f1",x"c2",x"86",x"cc"),
  1515 => (x"e9",x"49",x"bf",x"c0"),
  1516 => (x"9b",x"73",x"87",x"f5"),
  1517 => (x"c1",x"87",x"c8",x"02"),
  1518 => (x"c0",x"49",x"ee",x"e1"),
  1519 => (x"ff",x"87",x"fb",x"ef"),
  1520 => (x"1e",x"87",x"fa",x"df"),
  1521 => (x"48",x"d2",x"e2",x"c2"),
  1522 => (x"e3",x"c1",x"50",x"c0"),
  1523 => (x"c0",x"49",x"bf",x"d1"),
  1524 => (x"c0",x"87",x"c7",x"fe"),
  1525 => (x"1e",x"4f",x"26",x"48"),
  1526 => (x"c1",x"87",x"e5",x"c7"),
  1527 => (x"87",x"e5",x"fe",x"49"),
  1528 => (x"87",x"ce",x"eb",x"fe"),
  1529 => (x"cd",x"02",x"98",x"70"),
  1530 => (x"e9",x"f2",x"fe",x"87"),
  1531 => (x"02",x"98",x"70",x"87"),
  1532 => (x"4a",x"c1",x"87",x"c4"),
  1533 => (x"4a",x"c0",x"87",x"c2"),
  1534 => (x"ce",x"05",x"9a",x"72"),
  1535 => (x"c1",x"1e",x"c0",x"87"),
  1536 => (x"c0",x"49",x"eb",x"e0"),
  1537 => (x"c4",x"87",x"d1",x"fb"),
  1538 => (x"c1",x"87",x"fe",x"86"),
  1539 => (x"c0",x"87",x"ed",x"c2"),
  1540 => (x"f6",x"e0",x"c1",x"1e"),
  1541 => (x"ff",x"fa",x"c0",x"49"),
  1542 => (x"fe",x"1e",x"c0",x"87"),
  1543 => (x"49",x"70",x"87",x"e5"),
  1544 => (x"87",x"f4",x"fa",x"c0"),
  1545 => (x"f8",x"87",x"d8",x"c3"),
  1546 => (x"53",x"4f",x"26",x"8e"),
  1547 => (x"61",x"66",x"20",x"44"),
  1548 => (x"64",x"65",x"6c",x"69"),
  1549 => (x"6f",x"42",x"00",x"2e"),
  1550 => (x"6e",x"69",x"74",x"6f"),
  1551 => (x"2e",x"2e",x"2e",x"67"),
  1552 => (x"f2",x"c0",x"1e",x"00"),
  1553 => (x"87",x"fa",x"87",x"d5"),
  1554 => (x"c2",x"1e",x"4f",x"26"),
  1555 => (x"c0",x"48",x"c4",x"f1"),
  1556 => (x"c0",x"f1",x"c2",x"78"),
  1557 => (x"fd",x"78",x"c0",x"48"),
  1558 => (x"87",x"e5",x"87",x"fd"),
  1559 => (x"4f",x"26",x"48",x"c0"),
  1560 => (x"78",x"45",x"20",x"80"),
  1561 => (x"80",x"00",x"74",x"69"),
  1562 => (x"63",x"61",x"42",x"20"),
  1563 => (x"11",x"ff",x"00",x"6b"),
  1564 => (x"2c",x"59",x"00",x"00"),
  1565 => (x"00",x"00",x"00",x"00"),
  1566 => (x"00",x"11",x"ff",x"00"),
  1567 => (x"00",x"2c",x"77",x"00"),
  1568 => (x"00",x"00",x"00",x"00"),
  1569 => (x"00",x"00",x"11",x"ff"),
  1570 => (x"00",x"00",x"2c",x"95"),
  1571 => (x"ff",x"00",x"00",x"00"),
  1572 => (x"b3",x"00",x"00",x"11"),
  1573 => (x"00",x"00",x"00",x"2c"),
  1574 => (x"11",x"ff",x"00",x"00"),
  1575 => (x"2c",x"d1",x"00",x"00"),
  1576 => (x"00",x"00",x"00",x"00"),
  1577 => (x"00",x"11",x"ff",x"00"),
  1578 => (x"00",x"2c",x"ef",x"00"),
  1579 => (x"00",x"00",x"00",x"00"),
  1580 => (x"00",x"00",x"11",x"ff"),
  1581 => (x"00",x"00",x"2d",x"0d"),
  1582 => (x"ff",x"00",x"00",x"00"),
  1583 => (x"00",x"00",x"00",x"11"),
  1584 => (x"00",x"00",x"00",x"00"),
  1585 => (x"12",x"94",x"00",x"00"),
  1586 => (x"00",x"00",x"00",x"00"),
  1587 => (x"00",x"00",x"00",x"00"),
  1588 => (x"00",x"18",x"d5",x"00"),
  1589 => (x"4f",x"4f",x"42",x"00"),
  1590 => (x"20",x"20",x"20",x"54"),
  1591 => (x"4d",x"4f",x"52",x"20"),
  1592 => (x"61",x"6f",x"4c",x"00"),
  1593 => (x"2e",x"2a",x"20",x"64"),
  1594 => (x"f0",x"fe",x"1e",x"00"),
  1595 => (x"cd",x"78",x"c0",x"48"),
  1596 => (x"26",x"09",x"79",x"09"),
  1597 => (x"fe",x"1e",x"1e",x"4f"),
  1598 => (x"48",x"7e",x"bf",x"f0"),
  1599 => (x"1e",x"4f",x"26",x"26"),
  1600 => (x"c1",x"48",x"f0",x"fe"),
  1601 => (x"1e",x"4f",x"26",x"78"),
  1602 => (x"c0",x"48",x"f0",x"fe"),
  1603 => (x"1e",x"4f",x"26",x"78"),
  1604 => (x"52",x"c0",x"4a",x"71"),
  1605 => (x"0e",x"4f",x"26",x"52"),
  1606 => (x"5d",x"5c",x"5b",x"5e"),
  1607 => (x"71",x"86",x"f4",x"0e"),
  1608 => (x"7e",x"6d",x"97",x"4d"),
  1609 => (x"97",x"4c",x"a5",x"c1"),
  1610 => (x"a6",x"c8",x"48",x"6c"),
  1611 => (x"c4",x"48",x"6e",x"58"),
  1612 => (x"c5",x"05",x"a8",x"66"),
  1613 => (x"c0",x"48",x"ff",x"87"),
  1614 => (x"ca",x"ff",x"87",x"e6"),
  1615 => (x"49",x"a5",x"c2",x"87"),
  1616 => (x"71",x"4b",x"6c",x"97"),
  1617 => (x"6b",x"97",x"4b",x"a3"),
  1618 => (x"7e",x"6c",x"97",x"4b"),
  1619 => (x"80",x"c1",x"48",x"6e"),
  1620 => (x"c7",x"58",x"a6",x"c8"),
  1621 => (x"58",x"a6",x"cc",x"98"),
  1622 => (x"fe",x"7c",x"97",x"70"),
  1623 => (x"48",x"73",x"87",x"e1"),
  1624 => (x"4d",x"26",x"8e",x"f4"),
  1625 => (x"4b",x"26",x"4c",x"26"),
  1626 => (x"5e",x"0e",x"4f",x"26"),
  1627 => (x"f4",x"0e",x"5c",x"5b"),
  1628 => (x"d8",x"4c",x"71",x"86"),
  1629 => (x"ff",x"c3",x"4a",x"66"),
  1630 => (x"4b",x"a4",x"c2",x"9a"),
  1631 => (x"73",x"49",x"6c",x"97"),
  1632 => (x"51",x"72",x"49",x"a1"),
  1633 => (x"6e",x"7e",x"6c",x"97"),
  1634 => (x"c8",x"80",x"c1",x"48"),
  1635 => (x"98",x"c7",x"58",x"a6"),
  1636 => (x"70",x"58",x"a6",x"cc"),
  1637 => (x"ff",x"8e",x"f4",x"54"),
  1638 => (x"1e",x"1e",x"87",x"ca"),
  1639 => (x"e0",x"87",x"e8",x"fd"),
  1640 => (x"c0",x"49",x"4a",x"bf"),
  1641 => (x"02",x"99",x"c0",x"e0"),
  1642 => (x"1e",x"72",x"87",x"cb"),
  1643 => (x"49",x"eb",x"f4",x"c2"),
  1644 => (x"c4",x"87",x"f7",x"fe"),
  1645 => (x"87",x"fd",x"fc",x"86"),
  1646 => (x"c2",x"fd",x"7e",x"70"),
  1647 => (x"4f",x"26",x"26",x"87"),
  1648 => (x"eb",x"f4",x"c2",x"1e"),
  1649 => (x"87",x"c7",x"fd",x"49"),
  1650 => (x"49",x"da",x"e6",x"c1"),
  1651 => (x"c5",x"87",x"da",x"fc"),
  1652 => (x"4f",x"26",x"87",x"d9"),
  1653 => (x"5c",x"5b",x"5e",x"0e"),
  1654 => (x"f5",x"c2",x"0e",x"5d"),
  1655 => (x"c1",x"4a",x"bf",x"fe"),
  1656 => (x"49",x"bf",x"e8",x"e8"),
  1657 => (x"71",x"bc",x"72",x"4c"),
  1658 => (x"87",x"db",x"fc",x"4d"),
  1659 => (x"49",x"74",x"4b",x"c0"),
  1660 => (x"d5",x"02",x"99",x"d0"),
  1661 => (x"d0",x"49",x"75",x"87"),
  1662 => (x"c0",x"1e",x"71",x"99"),
  1663 => (x"fa",x"ee",x"c1",x"1e"),
  1664 => (x"12",x"82",x"73",x"4a"),
  1665 => (x"87",x"e4",x"c0",x"49"),
  1666 => (x"2c",x"c1",x"86",x"c8"),
  1667 => (x"ab",x"c8",x"83",x"2d"),
  1668 => (x"87",x"da",x"ff",x"04"),
  1669 => (x"c1",x"87",x"e8",x"fb"),
  1670 => (x"c2",x"48",x"e8",x"e8"),
  1671 => (x"78",x"bf",x"fe",x"f5"),
  1672 => (x"4c",x"26",x"4d",x"26"),
  1673 => (x"4f",x"26",x"4b",x"26"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"48",x"d0",x"ff",x"1e"),
  1676 => (x"ff",x"78",x"e1",x"c8"),
  1677 => (x"78",x"c5",x"48",x"d4"),
  1678 => (x"c3",x"02",x"66",x"c4"),
  1679 => (x"78",x"e0",x"c3",x"87"),
  1680 => (x"c6",x"02",x"66",x"c8"),
  1681 => (x"48",x"d4",x"ff",x"87"),
  1682 => (x"ff",x"78",x"f0",x"c3"),
  1683 => (x"78",x"71",x"48",x"d4"),
  1684 => (x"c8",x"48",x"d0",x"ff"),
  1685 => (x"e0",x"c0",x"78",x"e1"),
  1686 => (x"0e",x"4f",x"26",x"78"),
  1687 => (x"0e",x"5c",x"5b",x"5e"),
  1688 => (x"f4",x"c2",x"4c",x"71"),
  1689 => (x"ee",x"fa",x"49",x"eb"),
  1690 => (x"c0",x"4a",x"70",x"87"),
  1691 => (x"c2",x"04",x"aa",x"b7"),
  1692 => (x"e0",x"c3",x"87",x"e3"),
  1693 => (x"87",x"c9",x"05",x"aa"),
  1694 => (x"48",x"de",x"ec",x"c1"),
  1695 => (x"d4",x"c2",x"78",x"c1"),
  1696 => (x"aa",x"f0",x"c3",x"87"),
  1697 => (x"c1",x"87",x"c9",x"05"),
  1698 => (x"c1",x"48",x"da",x"ec"),
  1699 => (x"87",x"f5",x"c1",x"78"),
  1700 => (x"bf",x"de",x"ec",x"c1"),
  1701 => (x"72",x"87",x"c7",x"02"),
  1702 => (x"b3",x"c0",x"c2",x"4b"),
  1703 => (x"4b",x"72",x"87",x"c2"),
  1704 => (x"d1",x"05",x"9c",x"74"),
  1705 => (x"da",x"ec",x"c1",x"87"),
  1706 => (x"ec",x"c1",x"1e",x"bf"),
  1707 => (x"72",x"1e",x"bf",x"de"),
  1708 => (x"87",x"f8",x"fd",x"49"),
  1709 => (x"ec",x"c1",x"86",x"c8"),
  1710 => (x"c0",x"02",x"bf",x"da"),
  1711 => (x"49",x"73",x"87",x"e0"),
  1712 => (x"91",x"29",x"b7",x"c4"),
  1713 => (x"81",x"fa",x"ed",x"c1"),
  1714 => (x"9a",x"cf",x"4a",x"73"),
  1715 => (x"48",x"c1",x"92",x"c2"),
  1716 => (x"4a",x"70",x"30",x"72"),
  1717 => (x"48",x"72",x"ba",x"ff"),
  1718 => (x"79",x"70",x"98",x"69"),
  1719 => (x"49",x"73",x"87",x"db"),
  1720 => (x"91",x"29",x"b7",x"c4"),
  1721 => (x"81",x"fa",x"ed",x"c1"),
  1722 => (x"9a",x"cf",x"4a",x"73"),
  1723 => (x"48",x"c3",x"92",x"c2"),
  1724 => (x"4a",x"70",x"30",x"72"),
  1725 => (x"70",x"b0",x"69",x"48"),
  1726 => (x"de",x"ec",x"c1",x"79"),
  1727 => (x"c1",x"78",x"c0",x"48"),
  1728 => (x"c0",x"48",x"da",x"ec"),
  1729 => (x"eb",x"f4",x"c2",x"78"),
  1730 => (x"87",x"cb",x"f8",x"49"),
  1731 => (x"b7",x"c0",x"4a",x"70"),
  1732 => (x"dd",x"fd",x"03",x"aa"),
  1733 => (x"fc",x"48",x"c0",x"87"),
  1734 => (x"00",x"00",x"87",x"c8"),
  1735 => (x"00",x"00",x"00",x"00"),
  1736 => (x"71",x"1e",x"00",x"00"),
  1737 => (x"f2",x"fc",x"49",x"4a"),
  1738 => (x"1e",x"4f",x"26",x"87"),
  1739 => (x"49",x"72",x"4a",x"c0"),
  1740 => (x"ed",x"c1",x"91",x"c4"),
  1741 => (x"79",x"c0",x"81",x"fa"),
  1742 => (x"b7",x"d0",x"82",x"c1"),
  1743 => (x"87",x"ee",x"04",x"aa"),
  1744 => (x"5e",x"0e",x"4f",x"26"),
  1745 => (x"0e",x"5d",x"5c",x"5b"),
  1746 => (x"fa",x"f6",x"4d",x"71"),
  1747 => (x"c4",x"4a",x"75",x"87"),
  1748 => (x"c1",x"92",x"2a",x"b7"),
  1749 => (x"75",x"82",x"fa",x"ed"),
  1750 => (x"c2",x"9c",x"cf",x"4c"),
  1751 => (x"4b",x"49",x"6a",x"94"),
  1752 => (x"9b",x"c3",x"2b",x"74"),
  1753 => (x"30",x"74",x"48",x"c2"),
  1754 => (x"bc",x"ff",x"4c",x"70"),
  1755 => (x"98",x"71",x"48",x"74"),
  1756 => (x"ca",x"f6",x"7a",x"70"),
  1757 => (x"fa",x"48",x"73",x"87"),
  1758 => (x"00",x"00",x"87",x"e6"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"1e",x"16",x"00",x"00"),
  1775 => (x"36",x"2e",x"25",x"26"),
  1776 => (x"ff",x"1e",x"3e",x"3d"),
  1777 => (x"e1",x"c8",x"48",x"d0"),
  1778 => (x"ff",x"48",x"71",x"78"),
  1779 => (x"c4",x"78",x"08",x"d4"),
  1780 => (x"d4",x"ff",x"48",x"66"),
  1781 => (x"4f",x"26",x"78",x"08"),
  1782 => (x"c4",x"4a",x"71",x"1e"),
  1783 => (x"72",x"1e",x"49",x"66"),
  1784 => (x"87",x"de",x"ff",x"49"),
  1785 => (x"c0",x"48",x"d0",x"ff"),
  1786 => (x"26",x"26",x"78",x"e0"),
  1787 => (x"4a",x"71",x"1e",x"4f"),
  1788 => (x"c1",x"1e",x"66",x"c4"),
  1789 => (x"ff",x"49",x"a2",x"e0"),
  1790 => (x"66",x"c8",x"87",x"c8"),
  1791 => (x"29",x"b7",x"c8",x"49"),
  1792 => (x"71",x"48",x"d4",x"ff"),
  1793 => (x"48",x"d0",x"ff",x"78"),
  1794 => (x"26",x"78",x"e0",x"c0"),
  1795 => (x"ff",x"1e",x"4f",x"26"),
  1796 => (x"ff",x"c3",x"4a",x"d4"),
  1797 => (x"48",x"d0",x"ff",x"7a"),
  1798 => (x"de",x"78",x"e1",x"c8"),
  1799 => (x"f5",x"f4",x"c2",x"7a"),
  1800 => (x"48",x"49",x"7a",x"bf"),
  1801 => (x"7a",x"70",x"28",x"c8"),
  1802 => (x"28",x"d0",x"48",x"71"),
  1803 => (x"48",x"71",x"7a",x"70"),
  1804 => (x"7a",x"70",x"28",x"d8"),
  1805 => (x"c0",x"48",x"d0",x"ff"),
  1806 => (x"4f",x"26",x"78",x"e0"),
  1807 => (x"5c",x"5b",x"5e",x"0e"),
  1808 => (x"4c",x"71",x"0e",x"5d"),
  1809 => (x"bf",x"f5",x"f4",x"c2"),
  1810 => (x"2b",x"74",x"4b",x"4d"),
  1811 => (x"c1",x"9b",x"66",x"d0"),
  1812 => (x"ab",x"66",x"d4",x"83"),
  1813 => (x"c0",x"87",x"c2",x"04"),
  1814 => (x"d0",x"4a",x"74",x"4b"),
  1815 => (x"31",x"72",x"49",x"66"),
  1816 => (x"99",x"75",x"b9",x"ff"),
  1817 => (x"30",x"72",x"48",x"73"),
  1818 => (x"71",x"48",x"4a",x"70"),
  1819 => (x"f9",x"f4",x"c2",x"b0"),
  1820 => (x"87",x"da",x"fe",x"58"),
  1821 => (x"4c",x"26",x"4d",x"26"),
  1822 => (x"4f",x"26",x"4b",x"26"),
  1823 => (x"5c",x"5b",x"5e",x"0e"),
  1824 => (x"71",x"1e",x"0e",x"5d"),
  1825 => (x"f9",x"f4",x"c2",x"4c"),
  1826 => (x"c0",x"4a",x"c0",x"4b"),
  1827 => (x"d0",x"fe",x"49",x"f4"),
  1828 => (x"1e",x"74",x"87",x"f3"),
  1829 => (x"49",x"f9",x"f4",x"c2"),
  1830 => (x"87",x"c6",x"ed",x"fe"),
  1831 => (x"98",x"70",x"86",x"c4"),
  1832 => (x"87",x"ea",x"c0",x"02"),
  1833 => (x"4d",x"a6",x"1e",x"c4"),
  1834 => (x"f9",x"f4",x"c2",x"1e"),
  1835 => (x"f7",x"f2",x"fe",x"49"),
  1836 => (x"70",x"86",x"c8",x"87"),
  1837 => (x"87",x"d6",x"02",x"98"),
  1838 => (x"f4",x"c1",x"4a",x"75"),
  1839 => (x"4b",x"c4",x"49",x"c4"),
  1840 => (x"87",x"e6",x"ce",x"fe"),
  1841 => (x"ca",x"02",x"98",x"70"),
  1842 => (x"c0",x"48",x"c0",x"87"),
  1843 => (x"48",x"c0",x"87",x"ed"),
  1844 => (x"c0",x"87",x"e8",x"c0"),
  1845 => (x"c4",x"c1",x"87",x"f3"),
  1846 => (x"02",x"98",x"70",x"87"),
  1847 => (x"fc",x"c0",x"87",x"c8"),
  1848 => (x"05",x"98",x"70",x"87"),
  1849 => (x"f5",x"c2",x"87",x"f8"),
  1850 => (x"cc",x"02",x"bf",x"d9"),
  1851 => (x"f5",x"f4",x"c2",x"87"),
  1852 => (x"d9",x"f5",x"c2",x"48"),
  1853 => (x"d5",x"fc",x"78",x"bf"),
  1854 => (x"26",x"48",x"c1",x"87"),
  1855 => (x"4c",x"26",x"4d",x"26"),
  1856 => (x"4f",x"26",x"4b",x"26"),
  1857 => (x"43",x"52",x"41",x"5b"),
  1858 => (x"1e",x"c0",x"1e",x"00"),
  1859 => (x"49",x"f9",x"f4",x"c2"),
  1860 => (x"87",x"ed",x"ef",x"fe"),
  1861 => (x"48",x"d1",x"f5",x"c2"),
  1862 => (x"26",x"26",x"78",x"c0"),
  1863 => (x"5b",x"5e",x"0e",x"4f"),
  1864 => (x"f4",x"0e",x"5d",x"5c"),
  1865 => (x"48",x"a6",x"c4",x"86"),
  1866 => (x"f5",x"c2",x"78",x"c0"),
  1867 => (x"c3",x"48",x"bf",x"d1"),
  1868 => (x"d1",x"03",x"a8",x"b7"),
  1869 => (x"d1",x"f5",x"c2",x"87"),
  1870 => (x"80",x"c1",x"48",x"bf"),
  1871 => (x"58",x"d5",x"f5",x"c2"),
  1872 => (x"c6",x"48",x"fb",x"c0"),
  1873 => (x"f4",x"c2",x"87",x"e2"),
  1874 => (x"f4",x"fe",x"49",x"f9"),
  1875 => (x"4c",x"70",x"87",x"ee"),
  1876 => (x"bf",x"d1",x"f5",x"c2"),
  1877 => (x"02",x"8a",x"c3",x"4a"),
  1878 => (x"8a",x"c1",x"87",x"d8"),
  1879 => (x"87",x"cb",x"c5",x"02"),
  1880 => (x"f6",x"c2",x"02",x"8a"),
  1881 => (x"c1",x"02",x"8a",x"87"),
  1882 => (x"02",x"8a",x"87",x"cd"),
  1883 => (x"c5",x"87",x"e2",x"c3"),
  1884 => (x"4d",x"c0",x"87",x"e1"),
  1885 => (x"92",x"c4",x"4a",x"75"),
  1886 => (x"82",x"c6",x"fc",x"c1"),
  1887 => (x"48",x"cd",x"f5",x"c2"),
  1888 => (x"7e",x"70",x"80",x"75"),
  1889 => (x"4b",x"bf",x"97",x"6e"),
  1890 => (x"48",x"6e",x"4b",x"49"),
  1891 => (x"6a",x"50",x"a3",x"c1"),
  1892 => (x"cc",x"48",x"11",x"81"),
  1893 => (x"ac",x"70",x"58",x"a6"),
  1894 => (x"6e",x"87",x"c4",x"02"),
  1895 => (x"c8",x"50",x"c0",x"48"),
  1896 => (x"87",x"c7",x"05",x"66"),
  1897 => (x"48",x"d1",x"f5",x"c2"),
  1898 => (x"c1",x"78",x"a5",x"c4"),
  1899 => (x"ad",x"b7",x"c4",x"85"),
  1900 => (x"87",x"c0",x"ff",x"04"),
  1901 => (x"c2",x"87",x"dc",x"c4"),
  1902 => (x"48",x"bf",x"dd",x"f5"),
  1903 => (x"01",x"a8",x"b7",x"c8"),
  1904 => (x"ac",x"ca",x"87",x"d1"),
  1905 => (x"cd",x"87",x"cc",x"02"),
  1906 => (x"87",x"c7",x"02",x"ac"),
  1907 => (x"03",x"ac",x"b7",x"c0"),
  1908 => (x"c2",x"87",x"f3",x"c0"),
  1909 => (x"4b",x"bf",x"dd",x"f5"),
  1910 => (x"03",x"ab",x"b7",x"c8"),
  1911 => (x"f5",x"c2",x"87",x"d2"),
  1912 => (x"81",x"73",x"49",x"e1"),
  1913 => (x"c1",x"51",x"e0",x"c0"),
  1914 => (x"ab",x"b7",x"c8",x"83"),
  1915 => (x"87",x"ee",x"ff",x"04"),
  1916 => (x"48",x"e9",x"f5",x"c2"),
  1917 => (x"c1",x"50",x"d2",x"c1"),
  1918 => (x"cd",x"c1",x"50",x"cf"),
  1919 => (x"e4",x"50",x"c0",x"50"),
  1920 => (x"c3",x"78",x"c3",x"80"),
  1921 => (x"f5",x"c2",x"87",x"cd"),
  1922 => (x"48",x"49",x"bf",x"dd"),
  1923 => (x"f5",x"c2",x"80",x"c1"),
  1924 => (x"c4",x"48",x"58",x"e1"),
  1925 => (x"51",x"74",x"81",x"a0"),
  1926 => (x"c0",x"87",x"f8",x"c2"),
  1927 => (x"04",x"ac",x"b7",x"f0"),
  1928 => (x"f9",x"c0",x"87",x"da"),
  1929 => (x"d3",x"01",x"ac",x"b7"),
  1930 => (x"d5",x"f5",x"c2",x"87"),
  1931 => (x"91",x"ca",x"49",x"bf"),
  1932 => (x"f0",x"c0",x"4a",x"74"),
  1933 => (x"d5",x"f5",x"c2",x"8a"),
  1934 => (x"78",x"a1",x"72",x"48"),
  1935 => (x"c0",x"02",x"ac",x"ca"),
  1936 => (x"ac",x"cd",x"87",x"c6"),
  1937 => (x"87",x"cb",x"c2",x"05"),
  1938 => (x"48",x"d1",x"f5",x"c2"),
  1939 => (x"c2",x"c2",x"78",x"c3"),
  1940 => (x"b7",x"f0",x"c0",x"87"),
  1941 => (x"87",x"db",x"04",x"ac"),
  1942 => (x"ac",x"b7",x"f9",x"c0"),
  1943 => (x"87",x"d3",x"c0",x"01"),
  1944 => (x"bf",x"d9",x"f5",x"c2"),
  1945 => (x"74",x"91",x"d0",x"49"),
  1946 => (x"8a",x"f0",x"c0",x"4a"),
  1947 => (x"48",x"d9",x"f5",x"c2"),
  1948 => (x"c1",x"78",x"a1",x"72"),
  1949 => (x"04",x"ac",x"b7",x"c1"),
  1950 => (x"c1",x"87",x"db",x"c0"),
  1951 => (x"01",x"ac",x"b7",x"c6"),
  1952 => (x"c2",x"87",x"d3",x"c0"),
  1953 => (x"49",x"bf",x"d9",x"f5"),
  1954 => (x"4a",x"74",x"91",x"d0"),
  1955 => (x"c2",x"8a",x"f7",x"c0"),
  1956 => (x"72",x"48",x"d9",x"f5"),
  1957 => (x"ac",x"ca",x"78",x"a1"),
  1958 => (x"87",x"c6",x"c0",x"02"),
  1959 => (x"c0",x"05",x"ac",x"cd"),
  1960 => (x"f5",x"c2",x"87",x"f1"),
  1961 => (x"78",x"c3",x"48",x"d1"),
  1962 => (x"c0",x"87",x"e8",x"c0"),
  1963 => (x"c0",x"05",x"ac",x"e2"),
  1964 => (x"a6",x"c4",x"87",x"c9"),
  1965 => (x"78",x"fb",x"c0",x"48"),
  1966 => (x"ca",x"87",x"d8",x"c0"),
  1967 => (x"c6",x"c0",x"02",x"ac"),
  1968 => (x"05",x"ac",x"cd",x"87"),
  1969 => (x"c2",x"87",x"c9",x"c0"),
  1970 => (x"c3",x"48",x"d1",x"f5"),
  1971 => (x"87",x"c3",x"c0",x"78"),
  1972 => (x"c0",x"5c",x"a6",x"c8"),
  1973 => (x"c0",x"03",x"ac",x"b7"),
  1974 => (x"c0",x"48",x"87",x"c4"),
  1975 => (x"66",x"c4",x"87",x"ca"),
  1976 => (x"87",x"c6",x"f9",x"02"),
  1977 => (x"99",x"ff",x"c3",x"48"),
  1978 => (x"cf",x"f8",x"8e",x"f4"),
  1979 => (x"4e",x"4f",x"43",x"87"),
  1980 => (x"4d",x"00",x"3d",x"46"),
  1981 => (x"4e",x"00",x"44",x"4f"),
  1982 => (x"00",x"45",x"4d",x"41"),
  1983 => (x"41",x"46",x"45",x"44"),
  1984 => (x"3d",x"54",x"4c",x"55"),
  1985 => (x"1e",x"ed",x"00",x"30"),
  1986 => (x"1e",x"f3",x"00",x"00"),
  1987 => (x"1e",x"f7",x"00",x"00"),
  1988 => (x"1e",x"fc",x"00",x"00"),
  1989 => (x"ff",x"1e",x"00",x"00"),
  1990 => (x"c9",x"c8",x"48",x"d0"),
  1991 => (x"ff",x"48",x"71",x"78"),
  1992 => (x"26",x"78",x"08",x"d4"),
  1993 => (x"4a",x"71",x"1e",x"4f"),
  1994 => (x"ff",x"87",x"eb",x"49"),
  1995 => (x"78",x"c8",x"48",x"d0"),
  1996 => (x"73",x"1e",x"4f",x"26"),
  1997 => (x"c2",x"4b",x"71",x"1e"),
  1998 => (x"02",x"bf",x"f9",x"f5"),
  1999 => (x"eb",x"c2",x"87",x"c3"),
  2000 => (x"48",x"d0",x"ff",x"87"),
  2001 => (x"73",x"78",x"c9",x"c8"),
  2002 => (x"b1",x"e0",x"c0",x"49"),
  2003 => (x"71",x"48",x"d4",x"ff"),
  2004 => (x"ed",x"f5",x"c2",x"78"),
  2005 => (x"c8",x"78",x"c0",x"48"),
  2006 => (x"87",x"c5",x"02",x"66"),
  2007 => (x"c2",x"49",x"ff",x"c3"),
  2008 => (x"c2",x"49",x"c0",x"87"),
  2009 => (x"cc",x"59",x"f5",x"f5"),
  2010 => (x"87",x"c6",x"02",x"66"),
  2011 => (x"4a",x"d5",x"d5",x"c5"),
  2012 => (x"ff",x"cf",x"87",x"c4"),
  2013 => (x"f5",x"c2",x"4a",x"ff"),
  2014 => (x"f5",x"c2",x"5a",x"f9"),
  2015 => (x"78",x"c1",x"48",x"f9"),
  2016 => (x"4d",x"26",x"87",x"c4"),
  2017 => (x"4b",x"26",x"4c",x"26"),
  2018 => (x"5e",x"0e",x"4f",x"26"),
  2019 => (x"0e",x"5d",x"5c",x"5b"),
  2020 => (x"f5",x"c2",x"4a",x"71"),
  2021 => (x"72",x"4c",x"bf",x"f5"),
  2022 => (x"87",x"cb",x"02",x"9a"),
  2023 => (x"c1",x"91",x"c8",x"49"),
  2024 => (x"71",x"4b",x"e8",x"fc"),
  2025 => (x"c2",x"87",x"c4",x"83"),
  2026 => (x"c0",x"4b",x"e8",x"c0"),
  2027 => (x"74",x"49",x"13",x"4d"),
  2028 => (x"f1",x"f5",x"c2",x"99"),
  2029 => (x"d4",x"ff",x"b9",x"bf"),
  2030 => (x"c1",x"78",x"71",x"48"),
  2031 => (x"c8",x"85",x"2c",x"b7"),
  2032 => (x"e8",x"04",x"ad",x"b7"),
  2033 => (x"ed",x"f5",x"c2",x"87"),
  2034 => (x"80",x"c8",x"48",x"bf"),
  2035 => (x"58",x"f1",x"f5",x"c2"),
  2036 => (x"1e",x"87",x"ef",x"fe"),
  2037 => (x"4b",x"71",x"1e",x"73"),
  2038 => (x"02",x"9a",x"4a",x"13"),
  2039 => (x"49",x"72",x"87",x"cb"),
  2040 => (x"13",x"87",x"e7",x"fe"),
  2041 => (x"f5",x"05",x"9a",x"4a"),
  2042 => (x"87",x"da",x"fe",x"87"),
  2043 => (x"ed",x"f5",x"c2",x"1e"),
  2044 => (x"f5",x"c2",x"49",x"bf"),
  2045 => (x"a1",x"c1",x"48",x"ed"),
  2046 => (x"b7",x"c0",x"c4",x"78"),
  2047 => (x"87",x"db",x"03",x"a9"),
  2048 => (x"c2",x"48",x"d4",x"ff"),
  2049 => (x"78",x"bf",x"f1",x"f5"),
  2050 => (x"bf",x"ed",x"f5",x"c2"),
  2051 => (x"ed",x"f5",x"c2",x"49"),
  2052 => (x"78",x"a1",x"c1",x"48"),
  2053 => (x"a9",x"b7",x"c0",x"c4"),
  2054 => (x"ff",x"87",x"e5",x"04"),
  2055 => (x"78",x"c8",x"48",x"d0"),
  2056 => (x"48",x"f9",x"f5",x"c2"),
  2057 => (x"4f",x"26",x"78",x"c0"),
  2058 => (x"00",x"00",x"00",x"00"),
  2059 => (x"00",x"00",x"00",x"00"),
  2060 => (x"5f",x"00",x"00",x"00"),
  2061 => (x"00",x"00",x"00",x"5f"),
  2062 => (x"00",x"03",x"03",x"00"),
  2063 => (x"00",x"00",x"03",x"03"),
  2064 => (x"14",x"7f",x"7f",x"14"),
  2065 => (x"00",x"14",x"7f",x"7f"),
  2066 => (x"6b",x"2e",x"24",x"00"),
  2067 => (x"00",x"12",x"3a",x"6b"),
  2068 => (x"18",x"36",x"6a",x"4c"),
  2069 => (x"00",x"32",x"56",x"6c"),
  2070 => (x"59",x"4f",x"7e",x"30"),
  2071 => (x"40",x"68",x"3a",x"77"),
  2072 => (x"07",x"04",x"00",x"00"),
  2073 => (x"00",x"00",x"00",x"03"),
  2074 => (x"3e",x"1c",x"00",x"00"),
  2075 => (x"00",x"00",x"41",x"63"),
  2076 => (x"63",x"41",x"00",x"00"),
  2077 => (x"00",x"00",x"1c",x"3e"),
  2078 => (x"1c",x"3e",x"2a",x"08"),
  2079 => (x"08",x"2a",x"3e",x"1c"),
  2080 => (x"3e",x"08",x"08",x"00"),
  2081 => (x"00",x"08",x"08",x"3e"),
  2082 => (x"e0",x"80",x"00",x"00"),
  2083 => (x"00",x"00",x"00",x"60"),
  2084 => (x"08",x"08",x"08",x"00"),
  2085 => (x"00",x"08",x"08",x"08"),
  2086 => (x"60",x"00",x"00",x"00"),
  2087 => (x"00",x"00",x"00",x"60"),
  2088 => (x"18",x"30",x"60",x"40"),
  2089 => (x"01",x"03",x"06",x"0c"),
  2090 => (x"59",x"7f",x"3e",x"00"),
  2091 => (x"00",x"3e",x"7f",x"4d"),
  2092 => (x"7f",x"06",x"04",x"00"),
  2093 => (x"00",x"00",x"00",x"7f"),
  2094 => (x"71",x"63",x"42",x"00"),
  2095 => (x"00",x"46",x"4f",x"59"),
  2096 => (x"49",x"63",x"22",x"00"),
  2097 => (x"00",x"36",x"7f",x"49"),
  2098 => (x"13",x"16",x"1c",x"18"),
  2099 => (x"00",x"10",x"7f",x"7f"),
  2100 => (x"45",x"67",x"27",x"00"),
  2101 => (x"00",x"39",x"7d",x"45"),
  2102 => (x"4b",x"7e",x"3c",x"00"),
  2103 => (x"00",x"30",x"79",x"49"),
  2104 => (x"71",x"01",x"01",x"00"),
  2105 => (x"00",x"07",x"0f",x"79"),
  2106 => (x"49",x"7f",x"36",x"00"),
  2107 => (x"00",x"36",x"7f",x"49"),
  2108 => (x"49",x"4f",x"06",x"00"),
  2109 => (x"00",x"1e",x"3f",x"69"),
  2110 => (x"66",x"00",x"00",x"00"),
  2111 => (x"00",x"00",x"00",x"66"),
  2112 => (x"e6",x"80",x"00",x"00"),
  2113 => (x"00",x"00",x"00",x"66"),
  2114 => (x"14",x"08",x"08",x"00"),
  2115 => (x"00",x"22",x"22",x"14"),
  2116 => (x"14",x"14",x"14",x"00"),
  2117 => (x"00",x"14",x"14",x"14"),
  2118 => (x"14",x"22",x"22",x"00"),
  2119 => (x"00",x"08",x"08",x"14"),
  2120 => (x"51",x"03",x"02",x"00"),
  2121 => (x"00",x"06",x"0f",x"59"),
  2122 => (x"5d",x"41",x"7f",x"3e"),
  2123 => (x"00",x"1e",x"1f",x"55"),
  2124 => (x"09",x"7f",x"7e",x"00"),
  2125 => (x"00",x"7e",x"7f",x"09"),
  2126 => (x"49",x"7f",x"7f",x"00"),
  2127 => (x"00",x"36",x"7f",x"49"),
  2128 => (x"63",x"3e",x"1c",x"00"),
  2129 => (x"00",x"41",x"41",x"41"),
  2130 => (x"41",x"7f",x"7f",x"00"),
  2131 => (x"00",x"1c",x"3e",x"63"),
  2132 => (x"49",x"7f",x"7f",x"00"),
  2133 => (x"00",x"41",x"41",x"49"),
  2134 => (x"09",x"7f",x"7f",x"00"),
  2135 => (x"00",x"01",x"01",x"09"),
  2136 => (x"41",x"7f",x"3e",x"00"),
  2137 => (x"00",x"7a",x"7b",x"49"),
  2138 => (x"08",x"7f",x"7f",x"00"),
  2139 => (x"00",x"7f",x"7f",x"08"),
  2140 => (x"7f",x"41",x"00",x"00"),
  2141 => (x"00",x"00",x"41",x"7f"),
  2142 => (x"40",x"60",x"20",x"00"),
  2143 => (x"00",x"3f",x"7f",x"40"),
  2144 => (x"1c",x"08",x"7f",x"7f"),
  2145 => (x"00",x"41",x"63",x"36"),
  2146 => (x"40",x"7f",x"7f",x"00"),
  2147 => (x"00",x"40",x"40",x"40"),
  2148 => (x"0c",x"06",x"7f",x"7f"),
  2149 => (x"00",x"7f",x"7f",x"06"),
  2150 => (x"0c",x"06",x"7f",x"7f"),
  2151 => (x"00",x"7f",x"7f",x"18"),
  2152 => (x"41",x"7f",x"3e",x"00"),
  2153 => (x"00",x"3e",x"7f",x"41"),
  2154 => (x"09",x"7f",x"7f",x"00"),
  2155 => (x"00",x"06",x"0f",x"09"),
  2156 => (x"61",x"41",x"7f",x"3e"),
  2157 => (x"00",x"40",x"7e",x"7f"),
  2158 => (x"09",x"7f",x"7f",x"00"),
  2159 => (x"00",x"66",x"7f",x"19"),
  2160 => (x"4d",x"6f",x"26",x"00"),
  2161 => (x"00",x"32",x"7b",x"59"),
  2162 => (x"7f",x"01",x"01",x"00"),
  2163 => (x"00",x"01",x"01",x"7f"),
  2164 => (x"40",x"7f",x"3f",x"00"),
  2165 => (x"00",x"3f",x"7f",x"40"),
  2166 => (x"70",x"3f",x"0f",x"00"),
  2167 => (x"00",x"0f",x"3f",x"70"),
  2168 => (x"18",x"30",x"7f",x"7f"),
  2169 => (x"00",x"7f",x"7f",x"30"),
  2170 => (x"1c",x"36",x"63",x"41"),
  2171 => (x"41",x"63",x"36",x"1c"),
  2172 => (x"7c",x"06",x"03",x"01"),
  2173 => (x"01",x"03",x"06",x"7c"),
  2174 => (x"4d",x"59",x"71",x"61"),
  2175 => (x"00",x"41",x"43",x"47"),
  2176 => (x"7f",x"7f",x"00",x"00"),
  2177 => (x"00",x"00",x"41",x"41"),
  2178 => (x"0c",x"06",x"03",x"01"),
  2179 => (x"40",x"60",x"30",x"18"),
  2180 => (x"41",x"41",x"00",x"00"),
  2181 => (x"00",x"00",x"7f",x"7f"),
  2182 => (x"03",x"06",x"0c",x"08"),
  2183 => (x"00",x"08",x"0c",x"06"),
  2184 => (x"80",x"80",x"80",x"80"),
  2185 => (x"00",x"80",x"80",x"80"),
  2186 => (x"03",x"00",x"00",x"00"),
  2187 => (x"00",x"00",x"04",x"07"),
  2188 => (x"54",x"74",x"20",x"00"),
  2189 => (x"00",x"78",x"7c",x"54"),
  2190 => (x"44",x"7f",x"7f",x"00"),
  2191 => (x"00",x"38",x"7c",x"44"),
  2192 => (x"44",x"7c",x"38",x"00"),
  2193 => (x"00",x"00",x"44",x"44"),
  2194 => (x"44",x"7c",x"38",x"00"),
  2195 => (x"00",x"7f",x"7f",x"44"),
  2196 => (x"54",x"7c",x"38",x"00"),
  2197 => (x"00",x"18",x"5c",x"54"),
  2198 => (x"7f",x"7e",x"04",x"00"),
  2199 => (x"00",x"00",x"05",x"05"),
  2200 => (x"a4",x"bc",x"18",x"00"),
  2201 => (x"00",x"7c",x"fc",x"a4"),
  2202 => (x"04",x"7f",x"7f",x"00"),
  2203 => (x"00",x"78",x"7c",x"04"),
  2204 => (x"3d",x"00",x"00",x"00"),
  2205 => (x"00",x"00",x"40",x"7d"),
  2206 => (x"80",x"80",x"80",x"00"),
  2207 => (x"00",x"00",x"7d",x"fd"),
  2208 => (x"10",x"7f",x"7f",x"00"),
  2209 => (x"00",x"44",x"6c",x"38"),
  2210 => (x"3f",x"00",x"00",x"00"),
  2211 => (x"00",x"00",x"40",x"7f"),
  2212 => (x"18",x"0c",x"7c",x"7c"),
  2213 => (x"00",x"78",x"7c",x"0c"),
  2214 => (x"04",x"7c",x"7c",x"00"),
  2215 => (x"00",x"78",x"7c",x"04"),
  2216 => (x"44",x"7c",x"38",x"00"),
  2217 => (x"00",x"38",x"7c",x"44"),
  2218 => (x"24",x"fc",x"fc",x"00"),
  2219 => (x"00",x"18",x"3c",x"24"),
  2220 => (x"24",x"3c",x"18",x"00"),
  2221 => (x"00",x"fc",x"fc",x"24"),
  2222 => (x"04",x"7c",x"7c",x"00"),
  2223 => (x"00",x"08",x"0c",x"04"),
  2224 => (x"54",x"5c",x"48",x"00"),
  2225 => (x"00",x"20",x"74",x"54"),
  2226 => (x"7f",x"3f",x"04",x"00"),
  2227 => (x"00",x"00",x"44",x"44"),
  2228 => (x"40",x"7c",x"3c",x"00"),
  2229 => (x"00",x"7c",x"7c",x"40"),
  2230 => (x"60",x"3c",x"1c",x"00"),
  2231 => (x"00",x"1c",x"3c",x"60"),
  2232 => (x"30",x"60",x"7c",x"3c"),
  2233 => (x"00",x"3c",x"7c",x"60"),
  2234 => (x"10",x"38",x"6c",x"44"),
  2235 => (x"00",x"44",x"6c",x"38"),
  2236 => (x"e0",x"bc",x"1c",x"00"),
  2237 => (x"00",x"1c",x"3c",x"60"),
  2238 => (x"74",x"64",x"44",x"00"),
  2239 => (x"00",x"44",x"4c",x"5c"),
  2240 => (x"3e",x"08",x"08",x"00"),
  2241 => (x"00",x"41",x"41",x"77"),
  2242 => (x"7f",x"00",x"00",x"00"),
  2243 => (x"00",x"00",x"00",x"7f"),
  2244 => (x"77",x"41",x"41",x"00"),
  2245 => (x"00",x"08",x"08",x"3e"),
  2246 => (x"03",x"01",x"01",x"02"),
  2247 => (x"00",x"01",x"02",x"02"),
  2248 => (x"7f",x"7f",x"7f",x"7f"),
  2249 => (x"00",x"7f",x"7f",x"7f"),
  2250 => (x"1c",x"1c",x"08",x"08"),
  2251 => (x"7f",x"7f",x"3e",x"3e"),
  2252 => (x"3e",x"3e",x"7f",x"7f"),
  2253 => (x"08",x"08",x"1c",x"1c"),
  2254 => (x"7c",x"18",x"10",x"00"),
  2255 => (x"00",x"10",x"18",x"7c"),
  2256 => (x"7c",x"30",x"10",x"00"),
  2257 => (x"00",x"10",x"30",x"7c"),
  2258 => (x"60",x"60",x"30",x"10"),
  2259 => (x"00",x"06",x"1e",x"78"),
  2260 => (x"18",x"3c",x"66",x"42"),
  2261 => (x"00",x"42",x"66",x"3c"),
  2262 => (x"c2",x"6a",x"38",x"78"),
  2263 => (x"00",x"38",x"6c",x"c6"),
  2264 => (x"60",x"00",x"00",x"60"),
  2265 => (x"00",x"60",x"00",x"00"),
  2266 => (x"5c",x"5b",x"5e",x"0e"),
  2267 => (x"71",x"1e",x"0e",x"5d"),
  2268 => (x"ca",x"f6",x"c2",x"4c"),
  2269 => (x"4b",x"c0",x"4d",x"bf"),
  2270 => (x"ab",x"74",x"1e",x"c0"),
  2271 => (x"c4",x"87",x"c7",x"02"),
  2272 => (x"78",x"c0",x"48",x"a6"),
  2273 => (x"a6",x"c4",x"87",x"c5"),
  2274 => (x"c4",x"78",x"c1",x"48"),
  2275 => (x"49",x"73",x"1e",x"66"),
  2276 => (x"c8",x"87",x"df",x"ee"),
  2277 => (x"49",x"e0",x"c0",x"86"),
  2278 => (x"c4",x"87",x"ef",x"ef"),
  2279 => (x"49",x"6a",x"4a",x"a5"),
  2280 => (x"f1",x"87",x"f0",x"f0"),
  2281 => (x"85",x"cb",x"87",x"c6"),
  2282 => (x"b7",x"c8",x"83",x"c1"),
  2283 => (x"c7",x"ff",x"04",x"ab"),
  2284 => (x"4d",x"26",x"26",x"87"),
  2285 => (x"4b",x"26",x"4c",x"26"),
  2286 => (x"71",x"1e",x"4f",x"26"),
  2287 => (x"ce",x"f6",x"c2",x"4a"),
  2288 => (x"ce",x"f6",x"c2",x"5a"),
  2289 => (x"49",x"78",x"c7",x"48"),
  2290 => (x"26",x"87",x"dd",x"fe"),
  2291 => (x"1e",x"73",x"1e",x"4f"),
  2292 => (x"b7",x"c0",x"4a",x"71"),
  2293 => (x"87",x"d3",x"03",x"aa"),
  2294 => (x"bf",x"ed",x"dc",x"c2"),
  2295 => (x"c1",x"87",x"c4",x"05"),
  2296 => (x"c0",x"87",x"c2",x"4b"),
  2297 => (x"f1",x"dc",x"c2",x"4b"),
  2298 => (x"c2",x"87",x"c4",x"5b"),
  2299 => (x"c2",x"5a",x"f1",x"dc"),
  2300 => (x"4a",x"bf",x"ed",x"dc"),
  2301 => (x"c0",x"c1",x"9a",x"c1"),
  2302 => (x"e8",x"ec",x"49",x"a2"),
  2303 => (x"c2",x"48",x"fc",x"87"),
  2304 => (x"78",x"bf",x"ed",x"dc"),
  2305 => (x"1e",x"87",x"ef",x"fe"),
  2306 => (x"66",x"c4",x"4a",x"71"),
  2307 => (x"ff",x"49",x"72",x"1e"),
  2308 => (x"26",x"87",x"da",x"df"),
  2309 => (x"c2",x"1e",x"4f",x"26"),
  2310 => (x"49",x"bf",x"ed",x"dc"),
  2311 => (x"87",x"c2",x"dc",x"ff"),
  2312 => (x"48",x"c2",x"f6",x"c2"),
  2313 => (x"c2",x"78",x"bf",x"e8"),
  2314 => (x"ec",x"48",x"fe",x"f5"),
  2315 => (x"f6",x"c2",x"78",x"bf"),
  2316 => (x"49",x"4a",x"bf",x"c2"),
  2317 => (x"c8",x"99",x"ff",x"c3"),
  2318 => (x"48",x"72",x"2a",x"b7"),
  2319 => (x"f6",x"c2",x"b0",x"71"),
  2320 => (x"4f",x"26",x"58",x"ca"),
  2321 => (x"5c",x"5b",x"5e",x"0e"),
  2322 => (x"4b",x"71",x"0e",x"5d"),
  2323 => (x"c2",x"87",x"c7",x"ff"),
  2324 => (x"c0",x"48",x"fd",x"f5"),
  2325 => (x"ff",x"49",x"73",x"50"),
  2326 => (x"70",x"87",x"e7",x"db"),
  2327 => (x"9c",x"c2",x"4c",x"49"),
  2328 => (x"cb",x"49",x"ee",x"cb"),
  2329 => (x"49",x"70",x"87",x"cf"),
  2330 => (x"fd",x"f5",x"c2",x"4d"),
  2331 => (x"c1",x"05",x"bf",x"97"),
  2332 => (x"66",x"d0",x"87",x"e4"),
  2333 => (x"c6",x"f6",x"c2",x"49"),
  2334 => (x"d7",x"05",x"99",x"bf"),
  2335 => (x"49",x"66",x"d4",x"87"),
  2336 => (x"bf",x"fe",x"f5",x"c2"),
  2337 => (x"87",x"cc",x"05",x"99"),
  2338 => (x"da",x"ff",x"49",x"73"),
  2339 => (x"98",x"70",x"87",x"f4"),
  2340 => (x"87",x"c2",x"c1",x"02"),
  2341 => (x"fd",x"fd",x"4c",x"c1"),
  2342 => (x"ca",x"49",x"75",x"87"),
  2343 => (x"98",x"70",x"87",x"e3"),
  2344 => (x"c2",x"87",x"c6",x"02"),
  2345 => (x"c1",x"48",x"fd",x"f5"),
  2346 => (x"fd",x"f5",x"c2",x"50"),
  2347 => (x"c0",x"05",x"bf",x"97"),
  2348 => (x"f6",x"c2",x"87",x"e4"),
  2349 => (x"d0",x"49",x"bf",x"c6"),
  2350 => (x"ff",x"05",x"99",x"66"),
  2351 => (x"f5",x"c2",x"87",x"d6"),
  2352 => (x"d4",x"49",x"bf",x"fe"),
  2353 => (x"ff",x"05",x"99",x"66"),
  2354 => (x"49",x"73",x"87",x"ca"),
  2355 => (x"87",x"f2",x"d9",x"ff"),
  2356 => (x"fe",x"05",x"98",x"70"),
  2357 => (x"48",x"74",x"87",x"fe"),
  2358 => (x"0e",x"87",x"d7",x"fb"),
  2359 => (x"5d",x"5c",x"5b",x"5e"),
  2360 => (x"c0",x"86",x"f4",x"0e"),
  2361 => (x"bf",x"ec",x"4c",x"4d"),
  2362 => (x"48",x"a6",x"c4",x"7e"),
  2363 => (x"bf",x"ca",x"f6",x"c2"),
  2364 => (x"c0",x"1e",x"c1",x"78"),
  2365 => (x"fd",x"49",x"c7",x"1e"),
  2366 => (x"86",x"c8",x"87",x"ca"),
  2367 => (x"ce",x"02",x"98",x"70"),
  2368 => (x"fb",x"49",x"ff",x"87"),
  2369 => (x"da",x"c1",x"87",x"c7"),
  2370 => (x"f5",x"d8",x"ff",x"49"),
  2371 => (x"c2",x"4d",x"c1",x"87"),
  2372 => (x"bf",x"97",x"fd",x"f5"),
  2373 => (x"cd",x"87",x"c3",x"02"),
  2374 => (x"f6",x"c2",x"87",x"f9"),
  2375 => (x"c2",x"4b",x"bf",x"c2"),
  2376 => (x"05",x"bf",x"ed",x"dc"),
  2377 => (x"c3",x"87",x"eb",x"c0"),
  2378 => (x"d8",x"ff",x"49",x"fd"),
  2379 => (x"fa",x"c3",x"87",x"d4"),
  2380 => (x"cd",x"d8",x"ff",x"49"),
  2381 => (x"c3",x"49",x"73",x"87"),
  2382 => (x"1e",x"71",x"99",x"ff"),
  2383 => (x"c6",x"fb",x"49",x"c0"),
  2384 => (x"c8",x"49",x"73",x"87"),
  2385 => (x"1e",x"71",x"29",x"b7"),
  2386 => (x"fa",x"fa",x"49",x"c1"),
  2387 => (x"c6",x"86",x"c8",x"87"),
  2388 => (x"f6",x"c2",x"87",x"c1"),
  2389 => (x"9b",x"4b",x"bf",x"c6"),
  2390 => (x"c2",x"87",x"dd",x"02"),
  2391 => (x"49",x"bf",x"e9",x"dc"),
  2392 => (x"70",x"87",x"de",x"c7"),
  2393 => (x"87",x"c4",x"05",x"98"),
  2394 => (x"87",x"d2",x"4b",x"c0"),
  2395 => (x"c7",x"49",x"e0",x"c2"),
  2396 => (x"dc",x"c2",x"87",x"c3"),
  2397 => (x"87",x"c6",x"58",x"ed"),
  2398 => (x"48",x"e9",x"dc",x"c2"),
  2399 => (x"49",x"73",x"78",x"c0"),
  2400 => (x"ce",x"05",x"99",x"c2"),
  2401 => (x"49",x"eb",x"c3",x"87"),
  2402 => (x"87",x"f6",x"d6",x"ff"),
  2403 => (x"99",x"c2",x"49",x"70"),
  2404 => (x"fb",x"87",x"c2",x"02"),
  2405 => (x"c1",x"49",x"73",x"4c"),
  2406 => (x"87",x"ce",x"05",x"99"),
  2407 => (x"ff",x"49",x"f4",x"c3"),
  2408 => (x"70",x"87",x"df",x"d6"),
  2409 => (x"02",x"99",x"c2",x"49"),
  2410 => (x"4c",x"fa",x"87",x"c2"),
  2411 => (x"99",x"c8",x"49",x"73"),
  2412 => (x"c3",x"87",x"ce",x"05"),
  2413 => (x"d6",x"ff",x"49",x"f5"),
  2414 => (x"49",x"70",x"87",x"c8"),
  2415 => (x"d5",x"02",x"99",x"c2"),
  2416 => (x"ce",x"f6",x"c2",x"87"),
  2417 => (x"87",x"ca",x"02",x"bf"),
  2418 => (x"c2",x"88",x"c1",x"48"),
  2419 => (x"c0",x"58",x"d2",x"f6"),
  2420 => (x"4c",x"ff",x"87",x"c2"),
  2421 => (x"49",x"73",x"4d",x"c1"),
  2422 => (x"ce",x"05",x"99",x"c4"),
  2423 => (x"49",x"f2",x"c3",x"87"),
  2424 => (x"87",x"de",x"d5",x"ff"),
  2425 => (x"99",x"c2",x"49",x"70"),
  2426 => (x"c2",x"87",x"dc",x"02"),
  2427 => (x"7e",x"bf",x"ce",x"f6"),
  2428 => (x"a8",x"b7",x"c7",x"48"),
  2429 => (x"87",x"cb",x"c0",x"03"),
  2430 => (x"80",x"c1",x"48",x"6e"),
  2431 => (x"58",x"d2",x"f6",x"c2"),
  2432 => (x"fe",x"87",x"c2",x"c0"),
  2433 => (x"c3",x"4d",x"c1",x"4c"),
  2434 => (x"d4",x"ff",x"49",x"fd"),
  2435 => (x"49",x"70",x"87",x"f4"),
  2436 => (x"c0",x"02",x"99",x"c2"),
  2437 => (x"f6",x"c2",x"87",x"d5"),
  2438 => (x"c0",x"02",x"bf",x"ce"),
  2439 => (x"f6",x"c2",x"87",x"c9"),
  2440 => (x"78",x"c0",x"48",x"ce"),
  2441 => (x"fd",x"87",x"c2",x"c0"),
  2442 => (x"c3",x"4d",x"c1",x"4c"),
  2443 => (x"d4",x"ff",x"49",x"fa"),
  2444 => (x"49",x"70",x"87",x"d0"),
  2445 => (x"c0",x"02",x"99",x"c2"),
  2446 => (x"f6",x"c2",x"87",x"d9"),
  2447 => (x"c7",x"48",x"bf",x"ce"),
  2448 => (x"c0",x"03",x"a8",x"b7"),
  2449 => (x"f6",x"c2",x"87",x"c9"),
  2450 => (x"78",x"c7",x"48",x"ce"),
  2451 => (x"fc",x"87",x"c2",x"c0"),
  2452 => (x"c0",x"4d",x"c1",x"4c"),
  2453 => (x"c0",x"03",x"ac",x"b7"),
  2454 => (x"66",x"c4",x"87",x"d1"),
  2455 => (x"82",x"d8",x"c1",x"4a"),
  2456 => (x"c6",x"c0",x"02",x"6a"),
  2457 => (x"74",x"4b",x"6a",x"87"),
  2458 => (x"c0",x"0f",x"73",x"49"),
  2459 => (x"1e",x"f0",x"c3",x"1e"),
  2460 => (x"f7",x"49",x"da",x"c1"),
  2461 => (x"86",x"c8",x"87",x"ce"),
  2462 => (x"c0",x"02",x"98",x"70"),
  2463 => (x"a6",x"c8",x"87",x"e2"),
  2464 => (x"ce",x"f6",x"c2",x"48"),
  2465 => (x"66",x"c8",x"78",x"bf"),
  2466 => (x"c4",x"91",x"cb",x"49"),
  2467 => (x"80",x"71",x"48",x"66"),
  2468 => (x"bf",x"6e",x"7e",x"70"),
  2469 => (x"87",x"c8",x"c0",x"02"),
  2470 => (x"c8",x"4b",x"bf",x"6e"),
  2471 => (x"0f",x"73",x"49",x"66"),
  2472 => (x"c0",x"02",x"9d",x"75"),
  2473 => (x"f6",x"c2",x"87",x"c8"),
  2474 => (x"f2",x"49",x"bf",x"ce"),
  2475 => (x"dc",x"c2",x"87",x"fa"),
  2476 => (x"c0",x"02",x"bf",x"f1"),
  2477 => (x"c2",x"49",x"87",x"dd"),
  2478 => (x"98",x"70",x"87",x"c7"),
  2479 => (x"87",x"d3",x"c0",x"02"),
  2480 => (x"bf",x"ce",x"f6",x"c2"),
  2481 => (x"87",x"e0",x"f2",x"49"),
  2482 => (x"c0",x"f4",x"49",x"c0"),
  2483 => (x"f1",x"dc",x"c2",x"87"),
  2484 => (x"f4",x"78",x"c0",x"48"),
  2485 => (x"87",x"da",x"f3",x"8e"),
  2486 => (x"5c",x"5b",x"5e",x"0e"),
  2487 => (x"71",x"1e",x"0e",x"5d"),
  2488 => (x"ca",x"f6",x"c2",x"4c"),
  2489 => (x"cd",x"c1",x"49",x"bf"),
  2490 => (x"d1",x"c1",x"4d",x"a1"),
  2491 => (x"74",x"7e",x"69",x"81"),
  2492 => (x"87",x"cf",x"02",x"9c"),
  2493 => (x"74",x"4b",x"a5",x"c4"),
  2494 => (x"ca",x"f6",x"c2",x"7b"),
  2495 => (x"f9",x"f2",x"49",x"bf"),
  2496 => (x"74",x"7b",x"6e",x"87"),
  2497 => (x"87",x"c4",x"05",x"9c"),
  2498 => (x"87",x"c2",x"4b",x"c0"),
  2499 => (x"49",x"73",x"4b",x"c1"),
  2500 => (x"d4",x"87",x"fa",x"f2"),
  2501 => (x"87",x"c7",x"02",x"66"),
  2502 => (x"70",x"87",x"da",x"49"),
  2503 => (x"c0",x"87",x"c2",x"4a"),
  2504 => (x"f5",x"dc",x"c2",x"4a"),
  2505 => (x"c9",x"f2",x"26",x"5a"),
  2506 => (x"00",x"00",x"00",x"87"),
  2507 => (x"00",x"00",x"00",x"00"),
  2508 => (x"00",x"00",x"00",x"00"),
  2509 => (x"4a",x"71",x"1e",x"00"),
  2510 => (x"49",x"bf",x"c8",x"ff"),
  2511 => (x"26",x"48",x"a1",x"72"),
  2512 => (x"c8",x"ff",x"1e",x"4f"),
  2513 => (x"c0",x"fe",x"89",x"bf"),
  2514 => (x"c0",x"c0",x"c0",x"c0"),
  2515 => (x"87",x"c4",x"01",x"a9"),
  2516 => (x"87",x"c2",x"4a",x"c0"),
  2517 => (x"48",x"72",x"4a",x"c1"),
  2518 => (x"5e",x"0e",x"4f",x"26"),
  2519 => (x"0e",x"5d",x"5c",x"5b"),
  2520 => (x"ff",x"4d",x"71",x"1e"),
  2521 => (x"1e",x"75",x"4b",x"d4"),
  2522 => (x"49",x"d2",x"f6",x"c2"),
  2523 => (x"87",x"f2",x"c1",x"fe"),
  2524 => (x"7e",x"70",x"86",x"c4"),
  2525 => (x"ff",x"c3",x"02",x"6e"),
  2526 => (x"da",x"f6",x"c2",x"87"),
  2527 => (x"49",x"75",x"4c",x"bf"),
  2528 => (x"87",x"e0",x"db",x"fe"),
  2529 => (x"c0",x"05",x"a8",x"de"),
  2530 => (x"49",x"75",x"87",x"eb"),
  2531 => (x"87",x"ec",x"d3",x"ff"),
  2532 => (x"db",x"02",x"98",x"70"),
  2533 => (x"d5",x"f5",x"c2",x"87"),
  2534 => (x"e1",x"c0",x"1e",x"bf"),
  2535 => (x"f7",x"d0",x"ff",x"49"),
  2536 => (x"c2",x"86",x"c4",x"87"),
  2537 => (x"c0",x"48",x"d2",x"e2"),
  2538 => (x"e1",x"f5",x"c2",x"50"),
  2539 => (x"87",x"ea",x"fe",x"49"),
  2540 => (x"c5",x"c3",x"48",x"c1"),
  2541 => (x"48",x"d0",x"ff",x"87"),
  2542 => (x"c1",x"78",x"c5",x"c8"),
  2543 => (x"4a",x"c0",x"7b",x"d6"),
  2544 => (x"7b",x"bf",x"97",x"6e"),
  2545 => (x"80",x"c1",x"48",x"6e"),
  2546 => (x"82",x"c1",x"7e",x"70"),
  2547 => (x"aa",x"b7",x"e0",x"c0"),
  2548 => (x"87",x"ec",x"ff",x"04"),
  2549 => (x"c4",x"48",x"d0",x"ff"),
  2550 => (x"78",x"c5",x"c8",x"78"),
  2551 => (x"c1",x"7b",x"d3",x"c1"),
  2552 => (x"74",x"78",x"c4",x"7b"),
  2553 => (x"fd",x"c1",x"02",x"9c"),
  2554 => (x"ce",x"e4",x"c2",x"87"),
  2555 => (x"4d",x"c0",x"c8",x"7e"),
  2556 => (x"ac",x"b7",x"c0",x"8c"),
  2557 => (x"c8",x"87",x"c6",x"03"),
  2558 => (x"c0",x"4d",x"a4",x"c0"),
  2559 => (x"ff",x"f0",x"c2",x"4c"),
  2560 => (x"d0",x"49",x"bf",x"97"),
  2561 => (x"87",x"d2",x"02",x"99"),
  2562 => (x"f6",x"c2",x"1e",x"c0"),
  2563 => (x"c2",x"fe",x"49",x"d2"),
  2564 => (x"86",x"c4",x"87",x"ec"),
  2565 => (x"c0",x"4a",x"49",x"70"),
  2566 => (x"e4",x"c2",x"87",x"ef"),
  2567 => (x"f6",x"c2",x"1e",x"ce"),
  2568 => (x"c2",x"fe",x"49",x"d2"),
  2569 => (x"86",x"c4",x"87",x"d8"),
  2570 => (x"ff",x"4a",x"49",x"70"),
  2571 => (x"c5",x"c8",x"48",x"d0"),
  2572 => (x"7b",x"d4",x"c1",x"78"),
  2573 => (x"7b",x"bf",x"97",x"6e"),
  2574 => (x"80",x"c1",x"48",x"6e"),
  2575 => (x"8d",x"c1",x"7e",x"70"),
  2576 => (x"87",x"f0",x"ff",x"05"),
  2577 => (x"c4",x"48",x"d0",x"ff"),
  2578 => (x"05",x"9a",x"72",x"78"),
  2579 => (x"c0",x"87",x"c5",x"c0"),
  2580 => (x"87",x"e6",x"c0",x"48"),
  2581 => (x"f6",x"c2",x"1e",x"c1"),
  2582 => (x"ff",x"fd",x"49",x"d2"),
  2583 => (x"86",x"c4",x"87",x"ff"),
  2584 => (x"fe",x"05",x"9c",x"74"),
  2585 => (x"d0",x"ff",x"87",x"c3"),
  2586 => (x"78",x"c5",x"c8",x"48"),
  2587 => (x"c0",x"7b",x"d3",x"c1"),
  2588 => (x"c1",x"78",x"c4",x"7b"),
  2589 => (x"87",x"c2",x"c0",x"48"),
  2590 => (x"26",x"26",x"48",x"c0"),
  2591 => (x"26",x"4c",x"26",x"4d"),
  2592 => (x"1e",x"4f",x"26",x"4b"),
  2593 => (x"66",x"c4",x"4a",x"71"),
  2594 => (x"72",x"87",x"c5",x"05"),
  2595 => (x"87",x"ca",x"fb",x"49"),
  2596 => (x"1e",x"00",x"4f",x"26"),
  2597 => (x"bf",x"e1",x"e3",x"c2"),
  2598 => (x"c2",x"b9",x"c1",x"49"),
  2599 => (x"ff",x"59",x"e5",x"e3"),
  2600 => (x"ff",x"c3",x"48",x"d4"),
  2601 => (x"48",x"d0",x"ff",x"78"),
  2602 => (x"ff",x"78",x"e1",x"c8"),
  2603 => (x"78",x"c1",x"48",x"d4"),
  2604 => (x"78",x"71",x"31",x"c4"),
  2605 => (x"c0",x"48",x"d0",x"ff"),
  2606 => (x"4f",x"26",x"78",x"e0"),
  2607 => (x"d5",x"e3",x"c2",x"1e"),
  2608 => (x"d2",x"f6",x"c2",x"1e"),
  2609 => (x"d9",x"fc",x"fd",x"49"),
  2610 => (x"70",x"86",x"c4",x"87"),
  2611 => (x"87",x"c3",x"02",x"98"),
  2612 => (x"26",x"87",x"c0",x"ff"),
  2613 => (x"4b",x"35",x"31",x"4f"),
  2614 => (x"20",x"20",x"5a",x"48"),
  2615 => (x"47",x"46",x"43",x"20"),
  2616 => (x"00",x"00",x"00",x"00"),
  2617 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

