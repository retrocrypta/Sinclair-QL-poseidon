library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e8f6c287",
    12 => x"86c0c64e",
    13 => x"49e8f6c2",
    14 => x"48e8e3c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ffdf",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"ff1e4f26",
    53 => x"ffc348d4",
    54 => x"c4516878",
    55 => x"88c14866",
    56 => x"7058a6c8",
    57 => x"87eb0598",
    58 => x"731e4f26",
    59 => x"4bd4ff1e",
    60 => x"6b7bffc3",
    61 => x"7bffc34a",
    62 => x"32c8496b",
    63 => x"ffc3b172",
    64 => x"c84a6b7b",
    65 => x"c3b27131",
    66 => x"496b7bff",
    67 => x"b17232c8",
    68 => x"87c44871",
    69 => x"4c264d26",
    70 => x"4f264b26",
    71 => x"5c5b5e0e",
    72 => x"4a710e5d",
    73 => x"724cd4ff",
    74 => x"99ffc349",
    75 => x"e3c27c71",
    76 => x"c805bfe8",
    77 => x"4866d087",
    78 => x"a6d430c9",
    79 => x"4966d058",
    80 => x"ffc329d8",
    81 => x"d07c7199",
    82 => x"29d04966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"ffc329c8",
    86 => x"d07c7199",
    87 => x"ffc34966",
    88 => x"727c7199",
    89 => x"c329d049",
    90 => x"7c7199ff",
    91 => x"f0c94b6c",
    92 => x"ffc34dff",
    93 => x"87d005ab",
    94 => x"6c7cffc3",
    95 => x"028dc14b",
    96 => x"ffc387c6",
    97 => x"87f002ab",
    98 => x"c7fe4873",
    99 => x"49c01e87",
   100 => x"c348d4ff",
   101 => x"81c178ff",
   102 => x"a9b7c8c3",
   103 => x"2687f104",
   104 => x"1e731e4f",
   105 => x"f8c487e7",
   106 => x"1ec04bdf",
   107 => x"c1f0ffc0",
   108 => x"e7fd49f7",
   109 => x"c186c487",
   110 => x"eac005a8",
   111 => x"48d4ff87",
   112 => x"c178ffc3",
   113 => x"c0c0c0c0",
   114 => x"e1c01ec0",
   115 => x"49e9c1f0",
   116 => x"c487c9fd",
   117 => x"05987086",
   118 => x"d4ff87ca",
   119 => x"78ffc348",
   120 => x"87cb48c1",
   121 => x"c187e6fe",
   122 => x"fdfe058b",
   123 => x"fc48c087",
   124 => x"731e87e6",
   125 => x"48d4ff1e",
   126 => x"d378ffc3",
   127 => x"c01ec04b",
   128 => x"c1c1f0ff",
   129 => x"87d4fc49",
   130 => x"987086c4",
   131 => x"ff87ca05",
   132 => x"ffc348d4",
   133 => x"cb48c178",
   134 => x"87f1fd87",
   135 => x"ff058bc1",
   136 => x"48c087db",
   137 => x"0e87f1fb",
   138 => x"0e5c5b5e",
   139 => x"fd4cd4ff",
   140 => x"eac687db",
   141 => x"f0e1c01e",
   142 => x"fb49c8c1",
   143 => x"86c487de",
   144 => x"c802a8c1",
   145 => x"87eafe87",
   146 => x"e2c148c0",
   147 => x"87dafa87",
   148 => x"ffcf4970",
   149 => x"eac699ff",
   150 => x"87c802a9",
   151 => x"c087d3fe",
   152 => x"87cbc148",
   153 => x"c07cffc3",
   154 => x"f4fc4bf1",
   155 => x"02987087",
   156 => x"c087ebc0",
   157 => x"f0ffc01e",
   158 => x"fa49fac1",
   159 => x"86c487de",
   160 => x"d9059870",
   161 => x"7cffc387",
   162 => x"ffc3496c",
   163 => x"7c7c7c7c",
   164 => x"0299c0c1",
   165 => x"48c187c4",
   166 => x"48c087d5",
   167 => x"abc287d1",
   168 => x"c087c405",
   169 => x"c187c848",
   170 => x"fdfe058b",
   171 => x"f948c087",
   172 => x"731e87e4",
   173 => x"e8e3c21e",
   174 => x"c778c148",
   175 => x"48d0ff4b",
   176 => x"c8fb78c2",
   177 => x"48d0ff87",
   178 => x"1ec078c3",
   179 => x"c1d0e5c0",
   180 => x"c7f949c0",
   181 => x"c186c487",
   182 => x"87c105a8",
   183 => x"05abc24b",
   184 => x"48c087c5",
   185 => x"c187f9c0",
   186 => x"d0ff058b",
   187 => x"87f7fc87",
   188 => x"58ece3c2",
   189 => x"cd059870",
   190 => x"c01ec187",
   191 => x"d0c1f0ff",
   192 => x"87d8f849",
   193 => x"d4ff86c4",
   194 => x"78ffc348",
   195 => x"c287fec2",
   196 => x"ff58f0e3",
   197 => x"78c248d0",
   198 => x"c348d4ff",
   199 => x"48c178ff",
   200 => x"1e87f5f7",
   201 => x"ff4ad4ff",
   202 => x"d1c448d0",
   203 => x"7affc378",
   204 => x"f80589c1",
   205 => x"1e4f2687",
   206 => x"4b711e73",
   207 => x"dfcdeec5",
   208 => x"48d4ff4a",
   209 => x"6878ffc3",
   210 => x"a8fec348",
   211 => x"c187c502",
   212 => x"87ed058a",
   213 => x"c5059a72",
   214 => x"c048c087",
   215 => x"9b7387ea",
   216 => x"c887cc02",
   217 => x"49731e66",
   218 => x"c487e7f5",
   219 => x"c887c686",
   220 => x"eefe4966",
   221 => x"48d4ff87",
   222 => x"7878ffc3",
   223 => x"c5059b73",
   224 => x"48d0ff87",
   225 => x"48c178d0",
   226 => x"1e87cdf6",
   227 => x"4a711e73",
   228 => x"d4ff4bc0",
   229 => x"78ffc348",
   230 => x"c448d0ff",
   231 => x"d4ff78c3",
   232 => x"78ffc348",
   233 => x"ffc01e72",
   234 => x"49d1c1f0",
   235 => x"c487edf5",
   236 => x"05987086",
   237 => x"c0c887cd",
   238 => x"4966cc1e",
   239 => x"c487f8fd",
   240 => x"ff4b7086",
   241 => x"78c248d0",
   242 => x"cbf54873",
   243 => x"5b5e0e87",
   244 => x"c00e5d5c",
   245 => x"f0ffc01e",
   246 => x"f449c9c1",
   247 => x"1ed287fe",
   248 => x"49f0e3c2",
   249 => x"c887d0fd",
   250 => x"c14cc086",
   251 => x"acb7d284",
   252 => x"c287f804",
   253 => x"bf97f0e3",
   254 => x"99c0c349",
   255 => x"05a9c0c1",
   256 => x"c287e7c0",
   257 => x"bf97f7e3",
   258 => x"c231d049",
   259 => x"bf97f8e3",
   260 => x"7232c84a",
   261 => x"f9e3c2b1",
   262 => x"b14abf97",
   263 => x"ffcf4c71",
   264 => x"c19cffff",
   265 => x"c134ca84",
   266 => x"e3c287e7",
   267 => x"49bf97f9",
   268 => x"99c631c1",
   269 => x"97fae3c2",
   270 => x"b7c74abf",
   271 => x"c2b1722a",
   272 => x"bf97f5e3",
   273 => x"9dcf4d4a",
   274 => x"97f6e3c2",
   275 => x"9ac34abf",
   276 => x"e3c232ca",
   277 => x"4bbf97f7",
   278 => x"b27333c2",
   279 => x"97f8e3c2",
   280 => x"c0c34bbf",
   281 => x"2bb7c69b",
   282 => x"81c2b273",
   283 => x"307148c1",
   284 => x"48c14970",
   285 => x"4d703075",
   286 => x"84c14c72",
   287 => x"c0c89471",
   288 => x"cc06adb7",
   289 => x"b734c187",
   290 => x"b7c0c82d",
   291 => x"f4ff01ad",
   292 => x"f1487487",
   293 => x"5e0e87fe",
   294 => x"0e5d5c5b",
   295 => x"ecc286f8",
   296 => x"78c048d6",
   297 => x"1ecee4c2",
   298 => x"defb49c0",
   299 => x"7086c487",
   300 => x"87c50598",
   301 => x"cec948c0",
   302 => x"c14dc087",
   303 => x"caf5c07e",
   304 => x"e5c249bf",
   305 => x"c8714ac4",
   306 => x"87deee4b",
   307 => x"c2059870",
   308 => x"c07ec087",
   309 => x"49bfc6f5",
   310 => x"4ae0e5c2",
   311 => x"ee4bc871",
   312 => x"987087c8",
   313 => x"c087c205",
   314 => x"c0026e7e",
   315 => x"ebc287fd",
   316 => x"c24dbfd4",
   317 => x"bf9fccec",
   318 => x"d6c5487e",
   319 => x"c705a8ea",
   320 => x"d4ebc287",
   321 => x"87ce4dbf",
   322 => x"e9ca486e",
   323 => x"c502a8d5",
   324 => x"c748c087",
   325 => x"e4c287f1",
   326 => x"49751ece",
   327 => x"c487ecf9",
   328 => x"05987086",
   329 => x"48c087c5",
   330 => x"c087dcc7",
   331 => x"49bfc6f5",
   332 => x"4ae0e5c2",
   333 => x"ec4bc871",
   334 => x"987087f0",
   335 => x"c287c805",
   336 => x"c148d6ec",
   337 => x"c087da78",
   338 => x"49bfcaf5",
   339 => x"4ac4e5c2",
   340 => x"ec4bc871",
   341 => x"987087d4",
   342 => x"87c5c002",
   343 => x"e6c648c0",
   344 => x"ccecc287",
   345 => x"c149bf97",
   346 => x"c005a9d5",
   347 => x"ecc287cd",
   348 => x"49bf97cd",
   349 => x"02a9eac2",
   350 => x"c087c5c0",
   351 => x"87c7c648",
   352 => x"97cee4c2",
   353 => x"c3487ebf",
   354 => x"c002a8e9",
   355 => x"486e87ce",
   356 => x"02a8ebc3",
   357 => x"c087c5c0",
   358 => x"87ebc548",
   359 => x"97d9e4c2",
   360 => x"059949bf",
   361 => x"c287ccc0",
   362 => x"bf97dae4",
   363 => x"02a9c249",
   364 => x"c087c5c0",
   365 => x"87cfc548",
   366 => x"97dbe4c2",
   367 => x"ecc248bf",
   368 => x"4c7058d2",
   369 => x"c288c148",
   370 => x"c258d6ec",
   371 => x"bf97dce4",
   372 => x"c2817549",
   373 => x"bf97dde4",
   374 => x"7232c84a",
   375 => x"f0c27ea1",
   376 => x"786e48e3",
   377 => x"97dee4c2",
   378 => x"a6c848bf",
   379 => x"d6ecc258",
   380 => x"d4c202bf",
   381 => x"c6f5c087",
   382 => x"e5c249bf",
   383 => x"c8714ae0",
   384 => x"87e6e94b",
   385 => x"c0029870",
   386 => x"48c087c5",
   387 => x"c287f8c3",
   388 => x"4cbfceec",
   389 => x"5cf7f0c2",
   390 => x"97f3e4c2",
   391 => x"31c849bf",
   392 => x"97f2e4c2",
   393 => x"49a14abf",
   394 => x"97f4e4c2",
   395 => x"32d04abf",
   396 => x"c249a172",
   397 => x"bf97f5e4",
   398 => x"7232d84a",
   399 => x"66c449a1",
   400 => x"e3f0c291",
   401 => x"f0c281bf",
   402 => x"e4c259eb",
   403 => x"4abf97fb",
   404 => x"e4c232c8",
   405 => x"4bbf97fa",
   406 => x"e4c24aa2",
   407 => x"4bbf97fc",
   408 => x"a27333d0",
   409 => x"fde4c24a",
   410 => x"cf4bbf97",
   411 => x"7333d89b",
   412 => x"f0c24aa2",
   413 => x"f0c25aef",
   414 => x"c24abfeb",
   415 => x"c292748a",
   416 => x"7248eff0",
   417 => x"cac178a1",
   418 => x"e0e4c287",
   419 => x"c849bf97",
   420 => x"dfe4c231",
   421 => x"a14abf97",
   422 => x"deecc249",
   423 => x"daecc259",
   424 => x"31c549bf",
   425 => x"c981ffc7",
   426 => x"f7f0c229",
   427 => x"e5e4c259",
   428 => x"c84abf97",
   429 => x"e4e4c232",
   430 => x"a24bbf97",
   431 => x"9266c44a",
   432 => x"f0c2826e",
   433 => x"f0c25af3",
   434 => x"78c048eb",
   435 => x"48e7f0c2",
   436 => x"c278a172",
   437 => x"c248f7f0",
   438 => x"78bfebf0",
   439 => x"48fbf0c2",
   440 => x"bfeff0c2",
   441 => x"d6ecc278",
   442 => x"c9c002bf",
   443 => x"c4487487",
   444 => x"c07e7030",
   445 => x"f0c287c9",
   446 => x"c448bff3",
   447 => x"c27e7030",
   448 => x"6e48daec",
   449 => x"f848c178",
   450 => x"264d268e",
   451 => x"264b264c",
   452 => x"5b5e0e4f",
   453 => x"710e5d5c",
   454 => x"d6ecc24a",
   455 => x"87cb02bf",
   456 => x"2bc74b72",
   457 => x"ffc14c72",
   458 => x"7287c99c",
   459 => x"722bc84b",
   460 => x"9cffc34c",
   461 => x"bfe3f0c2",
   462 => x"c2f5c083",
   463 => x"d902abbf",
   464 => x"c6f5c087",
   465 => x"cee4c25b",
   466 => x"f049731e",
   467 => x"86c487fd",
   468 => x"c5059870",
   469 => x"c048c087",
   470 => x"ecc287e6",
   471 => x"d202bfd6",
   472 => x"c4497487",
   473 => x"cee4c291",
   474 => x"cf4d6981",
   475 => x"ffffffff",
   476 => x"7487cb9d",
   477 => x"c291c249",
   478 => x"9f81cee4",
   479 => x"48754d69",
   480 => x"0e87c6fe",
   481 => x"5d5c5b5e",
   482 => x"4d711e0e",
   483 => x"49c11ec0",
   484 => x"c487d7cf",
   485 => x"9c4c7086",
   486 => x"87c0c102",
   487 => x"4adeecc2",
   488 => x"eae24975",
   489 => x"02987087",
   490 => x"7487f1c0",
   491 => x"cb49754a",
   492 => x"87d0e34b",
   493 => x"c0029870",
   494 => x"1ec087e2",
   495 => x"c7029c74",
   496 => x"48a6c487",
   497 => x"87c578c0",
   498 => x"c148a6c4",
   499 => x"4966c478",
   500 => x"c487d7ce",
   501 => x"9c4c7086",
   502 => x"87c0ff05",
   503 => x"fc264874",
   504 => x"5e0e87e7",
   505 => x"0e5d5c5b",
   506 => x"9b4b711e",
   507 => x"c087c505",
   508 => x"87e5c148",
   509 => x"c04da3c8",
   510 => x"0266d47d",
   511 => x"66d487c7",
   512 => x"c505bf97",
   513 => x"c148c087",
   514 => x"66d487cf",
   515 => x"87f3fd49",
   516 => x"029c4c70",
   517 => x"dc87c0c1",
   518 => x"7d6949a4",
   519 => x"c449a4da",
   520 => x"699f4aa3",
   521 => x"d6ecc27a",
   522 => x"87d202bf",
   523 => x"9f49a4d4",
   524 => x"ffc04969",
   525 => x"487199ff",
   526 => x"7e7030d0",
   527 => x"7ec087c2",
   528 => x"6a48496e",
   529 => x"c07a7080",
   530 => x"49a3cc7b",
   531 => x"a3d0796a",
   532 => x"7479c049",
   533 => x"c087c248",
   534 => x"ecfa2648",
   535 => x"5b5e0e87",
   536 => x"710e5d5c",
   537 => x"c2f5c04c",
   538 => x"7478ff48",
   539 => x"cac1029c",
   540 => x"49a4c887",
   541 => x"c2c10269",
   542 => x"4a66d087",
   543 => x"d482496c",
   544 => x"66d05aa6",
   545 => x"ecc2b94d",
   546 => x"ff4abfd2",
   547 => x"719972ba",
   548 => x"e4c00299",
   549 => x"4ba4c487",
   550 => x"f4f9496b",
   551 => x"c27b7087",
   552 => x"49bfceec",
   553 => x"7c71816c",
   554 => x"ecc2b975",
   555 => x"ff4abfd2",
   556 => x"719972ba",
   557 => x"dcff0599",
   558 => x"f97c7587",
   559 => x"731e87cb",
   560 => x"9b4b711e",
   561 => x"c887c702",
   562 => x"056949a3",
   563 => x"48c087c5",
   564 => x"c287ebc0",
   565 => x"4abfe7f0",
   566 => x"6949a3c4",
   567 => x"c289c249",
   568 => x"91bfceec",
   569 => x"c24aa271",
   570 => x"49bfd2ec",
   571 => x"a271996b",
   572 => x"1e66c84a",
   573 => x"d2ea4972",
   574 => x"7086c487",
   575 => x"ccf84849",
   576 => x"5b5e0e87",
   577 => x"1e0e5d5c",
   578 => x"66d44b71",
   579 => x"732cc94c",
   580 => x"cfc1029b",
   581 => x"49a3c887",
   582 => x"c7c10269",
   583 => x"4da3d087",
   584 => x"c27d66d4",
   585 => x"49bfd2ec",
   586 => x"4a6bb9ff",
   587 => x"ac717e99",
   588 => x"c087cd03",
   589 => x"a3cc7d7b",
   590 => x"49a3c44a",
   591 => x"87c2796a",
   592 => x"9c748c72",
   593 => x"4987dd02",
   594 => x"fc49731e",
   595 => x"86c487cf",
   596 => x"c74966d4",
   597 => x"cb0299ff",
   598 => x"cee4c287",
   599 => x"fd49731e",
   600 => x"86c487dc",
   601 => x"87e1f626",
   602 => x"5c5b5e0e",
   603 => x"86f00e5d",
   604 => x"c059a6d0",
   605 => x"cc4b66e4",
   606 => x"87ca0266",
   607 => x"7080c848",
   608 => x"05bf6e7e",
   609 => x"48c087c5",
   610 => x"cc87ecc3",
   611 => x"84d04c66",
   612 => x"a6c44973",
   613 => x"c4786c48",
   614 => x"80c48166",
   615 => x"c878bf6e",
   616 => x"c606a966",
   617 => x"66c44987",
   618 => x"c04b7189",
   619 => x"c401abb7",
   620 => x"c2c34887",
   621 => x"4866c487",
   622 => x"7098ffc7",
   623 => x"c1026e7e",
   624 => x"c0c887c9",
   625 => x"71896e49",
   626 => x"cee4c24a",
   627 => x"73856e4d",
   628 => x"c106aab7",
   629 => x"49724a87",
   630 => x"8066c448",
   631 => x"8b727c70",
   632 => x"718ac149",
   633 => x"87d90299",
   634 => x"4866e0c0",
   635 => x"e0c05015",
   636 => x"80c14866",
   637 => x"58a6e4c0",
   638 => x"8ac14972",
   639 => x"e7059971",
   640 => x"d01ec187",
   641 => x"d4f94966",
   642 => x"c086c487",
   643 => x"c106abb7",
   644 => x"e0c087e3",
   645 => x"ffc74d66",
   646 => x"c006abb7",
   647 => x"1e7587e2",
   648 => x"fa4966d0",
   649 => x"c0c887d8",
   650 => x"c8486c85",
   651 => x"7c7080c0",
   652 => x"c18bc0c8",
   653 => x"4966d41e",
   654 => x"c887e2f8",
   655 => x"87eec086",
   656 => x"1ecee4c2",
   657 => x"f94966d0",
   658 => x"86c487f4",
   659 => x"4acee4c2",
   660 => x"6c484973",
   661 => x"737c7080",
   662 => x"718bc149",
   663 => x"87ce0299",
   664 => x"c17d9712",
   665 => x"c1497385",
   666 => x"0599718b",
   667 => x"b7c087f2",
   668 => x"e1fe01ab",
   669 => x"f048c187",
   670 => x"87cdf28e",
   671 => x"5c5b5e0e",
   672 => x"4b710e5d",
   673 => x"87c7029b",
   674 => x"6d4da3c8",
   675 => x"ff87c505",
   676 => x"87fdc048",
   677 => x"6c4ca3d0",
   678 => x"99ffc749",
   679 => x"6c87d805",
   680 => x"c187c902",
   681 => x"f649731e",
   682 => x"86c487f3",
   683 => x"1ecee4c2",
   684 => x"c9f84973",
   685 => x"6c86c487",
   686 => x"04aa6d4a",
   687 => x"48ff87c4",
   688 => x"a2c187cf",
   689 => x"c749727c",
   690 => x"e4c299ff",
   691 => x"699781ce",
   692 => x"87f5f048",
   693 => x"711e731e",
   694 => x"c0029b4b",
   695 => x"f0c287e4",
   696 => x"4a735bfb",
   697 => x"ecc28ac2",
   698 => x"9249bfce",
   699 => x"bfe7f0c2",
   700 => x"c2807248",
   701 => x"7158fff0",
   702 => x"c230c448",
   703 => x"c058deec",
   704 => x"f0c287ed",
   705 => x"f0c248f7",
   706 => x"c278bfeb",
   707 => x"c248fbf0",
   708 => x"78bfeff0",
   709 => x"bfd6ecc2",
   710 => x"c287c902",
   711 => x"49bfceec",
   712 => x"87c731c4",
   713 => x"bff3f0c2",
   714 => x"c231c449",
   715 => x"ef59deec",
   716 => x"5e0e87db",
   717 => x"710e5c5b",
   718 => x"724bc04a",
   719 => x"e1c0029a",
   720 => x"49a2da87",
   721 => x"c24b699f",
   722 => x"02bfd6ec",
   723 => x"a2d487cf",
   724 => x"49699f49",
   725 => x"ffffc04c",
   726 => x"c234d09c",
   727 => x"744cc087",
   728 => x"4973b349",
   729 => x"ee87edfd",
   730 => x"5e0e87e1",
   731 => x"0e5d5c5b",
   732 => x"4a7186f4",
   733 => x"9a727ec0",
   734 => x"c287d802",
   735 => x"c048cae4",
   736 => x"c2e4c278",
   737 => x"fbf0c248",
   738 => x"e4c278bf",
   739 => x"f0c248c6",
   740 => x"c278bff7",
   741 => x"c048ebec",
   742 => x"daecc250",
   743 => x"e4c249bf",
   744 => x"714abfca",
   745 => x"c0c403aa",
   746 => x"cf497287",
   747 => x"e1c00599",
   748 => x"cee4c287",
   749 => x"c2e4c21e",
   750 => x"e4c249bf",
   751 => x"a1c148c2",
   752 => x"dfff7178",
   753 => x"86c487c5",
   754 => x"48fef4c0",
   755 => x"78cee4c2",
   756 => x"f4c087cc",
   757 => x"c048bffe",
   758 => x"f5c080e0",
   759 => x"e4c258c2",
   760 => x"c148bfca",
   761 => x"cee4c280",
   762 => x"0d3e2758",
   763 => x"97bf0000",
   764 => x"029d4dbf",
   765 => x"c387e2c2",
   766 => x"c202ade5",
   767 => x"f4c087db",
   768 => x"cb4bbffe",
   769 => x"4c1149a3",
   770 => x"c105accf",
   771 => x"497587d2",
   772 => x"89c199df",
   773 => x"ecc291cd",
   774 => x"a3c181de",
   775 => x"c351124a",
   776 => x"51124aa3",
   777 => x"124aa3c5",
   778 => x"4aa3c751",
   779 => x"a3c95112",
   780 => x"ce51124a",
   781 => x"51124aa3",
   782 => x"124aa3d0",
   783 => x"4aa3d251",
   784 => x"a3d45112",
   785 => x"d651124a",
   786 => x"51124aa3",
   787 => x"124aa3d8",
   788 => x"4aa3dc51",
   789 => x"a3de5112",
   790 => x"c151124a",
   791 => x"87f9c07e",
   792 => x"99c84974",
   793 => x"87eac005",
   794 => x"99d04974",
   795 => x"dc87d005",
   796 => x"cac00266",
   797 => x"dc497387",
   798 => x"98700f66",
   799 => x"6e87d302",
   800 => x"87c6c005",
   801 => x"48deecc2",
   802 => x"f4c050c0",
   803 => x"c248bffe",
   804 => x"ecc287e7",
   805 => x"50c048eb",
   806 => x"daecc27e",
   807 => x"e4c249bf",
   808 => x"714abfca",
   809 => x"c0fc04aa",
   810 => x"fbf0c287",
   811 => x"c8c005bf",
   812 => x"d6ecc287",
   813 => x"fec102bf",
   814 => x"c2f5c087",
   815 => x"c278ff48",
   816 => x"49bfc6e4",
   817 => x"7087cae9",
   818 => x"cae4c249",
   819 => x"48a6c459",
   820 => x"bfc6e4c2",
   821 => x"d6ecc278",
   822 => x"d8c002bf",
   823 => x"4966c487",
   824 => x"ffffffcf",
   825 => x"02a999f8",
   826 => x"c087c5c0",
   827 => x"87e1c04d",
   828 => x"dcc04dc1",
   829 => x"4966c487",
   830 => x"99f8ffcf",
   831 => x"c8c002a9",
   832 => x"48a6c887",
   833 => x"c5c078c0",
   834 => x"48a6c887",
   835 => x"66c878c1",
   836 => x"059d754d",
   837 => x"c487e0c0",
   838 => x"89c24966",
   839 => x"bfceecc2",
   840 => x"f0c2914a",
   841 => x"c24abfe7",
   842 => x"7248c2e4",
   843 => x"e4c278a1",
   844 => x"78c048ca",
   845 => x"c087e2f9",
   846 => x"e78ef448",
   847 => x"000087cb",
   848 => x"ffff0000",
   849 => x"0d4effff",
   850 => x"0d570000",
   851 => x"41460000",
   852 => x"20323354",
   853 => x"46002020",
   854 => x"36315441",
   855 => x"00202020",
   856 => x"c0f1c21e",
   857 => x"a8dd48bf",
   858 => x"c087c905",
   859 => x"7087eefe",
   860 => x"87c84a49",
   861 => x"c348d4ff",
   862 => x"4a6878ff",
   863 => x"4f264872",
   864 => x"c0f1c21e",
   865 => x"a8dd48bf",
   866 => x"c087c605",
   867 => x"d987fafd",
   868 => x"48d4ff87",
   869 => x"ff78ffc3",
   870 => x"e1c848d0",
   871 => x"48d4ff78",
   872 => x"f0c278d4",
   873 => x"d4ff48ff",
   874 => x"4f2650bf",
   875 => x"48d0ff1e",
   876 => x"2678e0c0",
   877 => x"e7fe1e4f",
   878 => x"99497087",
   879 => x"c087c602",
   880 => x"f105a9fb",
   881 => x"26487187",
   882 => x"5b5e0e4f",
   883 => x"4b710e5c",
   884 => x"cbfe4cc0",
   885 => x"99497087",
   886 => x"87f9c002",
   887 => x"02a9ecc0",
   888 => x"c087f2c0",
   889 => x"c002a9fb",
   890 => x"66cc87eb",
   891 => x"c703acb7",
   892 => x"0266d087",
   893 => x"537187c2",
   894 => x"c2029971",
   895 => x"fd84c187",
   896 => x"497087de",
   897 => x"87cd0299",
   898 => x"02a9ecc0",
   899 => x"fbc087c7",
   900 => x"d5ff05a9",
   901 => x"0266d087",
   902 => x"97c087c3",
   903 => x"a9ecc07b",
   904 => x"7487c405",
   905 => x"7487c54a",
   906 => x"8a0ac04a",
   907 => x"87c24872",
   908 => x"4c264d26",
   909 => x"4f264b26",
   910 => x"87e4fc1e",
   911 => x"f0c04970",
   912 => x"ca04a9b7",
   913 => x"b7f9c087",
   914 => x"87c301a9",
   915 => x"c189f0c0",
   916 => x"04a9b7c1",
   917 => x"dac187ca",
   918 => x"c301a9b7",
   919 => x"89f7c087",
   920 => x"4f264871",
   921 => x"5c5b5e0e",
   922 => x"ff4a710e",
   923 => x"49724cd4",
   924 => x"7087eac0",
   925 => x"c2029b4b",
   926 => x"ff8bc187",
   927 => x"c5c848d0",
   928 => x"7cd5c178",
   929 => x"31c64973",
   930 => x"97d2e2c2",
   931 => x"71484abf",
   932 => x"ff7c70b0",
   933 => x"78c448d0",
   934 => x"d5fe4873",
   935 => x"5b5e0e87",
   936 => x"f40e5d5c",
   937 => x"c44c7186",
   938 => x"78c048a6",
   939 => x"6e7ea4c8",
   940 => x"c149bf97",
   941 => x"dd05a9c1",
   942 => x"49a4c987",
   943 => x"c1496997",
   944 => x"d105a9d2",
   945 => x"49a4ca87",
   946 => x"c1496997",
   947 => x"c505a9c3",
   948 => x"c248df87",
   949 => x"e7fa87e1",
   950 => x"c04bc087",
   951 => x"bf97fcfd",
   952 => x"04a9c049",
   953 => x"ccfb87cf",
   954 => x"c083c187",
   955 => x"bf97fcfd",
   956 => x"f106ab49",
   957 => x"fcfdc087",
   958 => x"cf02bf97",
   959 => x"87e0f987",
   960 => x"02994970",
   961 => x"ecc087c6",
   962 => x"87f105a9",
   963 => x"cff94bc0",
   964 => x"f94d7087",
   965 => x"a6cc87ca",
   966 => x"87c4f958",
   967 => x"83c14a70",
   968 => x"49bf976e",
   969 => x"87c702ad",
   970 => x"05adffc0",
   971 => x"c987eac0",
   972 => x"699749a4",
   973 => x"a966c849",
   974 => x"4887c702",
   975 => x"05a8ffc0",
   976 => x"a4ca87d7",
   977 => x"49699749",
   978 => x"87c602aa",
   979 => x"05aaffc0",
   980 => x"a6c487c7",
   981 => x"d378c148",
   982 => x"adecc087",
   983 => x"c087c602",
   984 => x"c705adfb",
   985 => x"c44bc087",
   986 => x"78c148a6",
   987 => x"fe0266c4",
   988 => x"f7f887dc",
   989 => x"f4487387",
   990 => x"87f4fa8e",
   991 => x"5b5e0e00",
   992 => x"1e0e5d5c",
   993 => x"4cc04b71",
   994 => x"c004ab4d",
   995 => x"fac087e8",
   996 => x"9d751edd",
   997 => x"c087c402",
   998 => x"c187c24a",
   999 => x"ef49724a",
  1000 => x"86c487c8",
  1001 => x"84c17e70",
  1002 => x"87c2056e",
  1003 => x"85c14c73",
  1004 => x"ff06ac73",
  1005 => x"486e87d8",
  1006 => x"264d2626",
  1007 => x"264b264c",
  1008 => x"5b5e0e4f",
  1009 => x"1e0e5d5c",
  1010 => x"de494c71",
  1011 => x"d9f1c291",
  1012 => x"9785714d",
  1013 => x"ddc1026d",
  1014 => x"c4f1c287",
  1015 => x"82744abf",
  1016 => x"d8fe4972",
  1017 => x"6e7e7087",
  1018 => x"87f3c002",
  1019 => x"4bccf1c2",
  1020 => x"49cb4a6e",
  1021 => x"87f0c2ff",
  1022 => x"93cb4b74",
  1023 => x"83eee1c1",
  1024 => x"c0c183c4",
  1025 => x"49747bfa",
  1026 => x"87dccdc1",
  1027 => x"f1c27b75",
  1028 => x"49bf97d8",
  1029 => x"ccf1c21e",
  1030 => x"e6e1c149",
  1031 => x"7486c487",
  1032 => x"c3cdc149",
  1033 => x"c149c087",
  1034 => x"c287e2ce",
  1035 => x"c048c0f1",
  1036 => x"dd49c178",
  1037 => x"fd2687cf",
  1038 => x"6f4c87ff",
  1039 => x"6e696461",
  1040 => x"2e2e2e67",
  1041 => x"5b5e0e00",
  1042 => x"4b710e5c",
  1043 => x"c4f1c24a",
  1044 => x"497282bf",
  1045 => x"7087e6fc",
  1046 => x"c4029c4c",
  1047 => x"d1eb4987",
  1048 => x"c4f1c287",
  1049 => x"c178c048",
  1050 => x"87d9dc49",
  1051 => x"0e87ccfd",
  1052 => x"5d5c5b5e",
  1053 => x"c286f40e",
  1054 => x"c04dcee4",
  1055 => x"48a6c44c",
  1056 => x"f1c278c0",
  1057 => x"c049bfc4",
  1058 => x"c1c106a9",
  1059 => x"cee4c287",
  1060 => x"c0029848",
  1061 => x"fac087f8",
  1062 => x"66c81edd",
  1063 => x"c487c702",
  1064 => x"78c048a6",
  1065 => x"a6c487c5",
  1066 => x"c478c148",
  1067 => x"f9ea4966",
  1068 => x"7086c487",
  1069 => x"c484c14d",
  1070 => x"80c14866",
  1071 => x"c258a6c8",
  1072 => x"49bfc4f1",
  1073 => x"87c603ac",
  1074 => x"ff059d75",
  1075 => x"4cc087c8",
  1076 => x"c3029d75",
  1077 => x"fac087e0",
  1078 => x"66c81edd",
  1079 => x"cc87c702",
  1080 => x"78c048a6",
  1081 => x"a6cc87c5",
  1082 => x"cc78c148",
  1083 => x"f9e94966",
  1084 => x"7086c487",
  1085 => x"c2026e7e",
  1086 => x"496e87e9",
  1087 => x"699781cb",
  1088 => x"0299d049",
  1089 => x"c187d6c1",
  1090 => x"744ac5c1",
  1091 => x"c191cb49",
  1092 => x"7281eee1",
  1093 => x"c381c879",
  1094 => x"497451ff",
  1095 => x"f1c291de",
  1096 => x"85714dd9",
  1097 => x"7d97c1c2",
  1098 => x"c049a5c1",
  1099 => x"ecc251e0",
  1100 => x"02bf97de",
  1101 => x"84c187d2",
  1102 => x"c24ba5c2",
  1103 => x"db4adeec",
  1104 => x"e3fdfe49",
  1105 => x"87dbc187",
  1106 => x"c049a5cd",
  1107 => x"c284c151",
  1108 => x"4a6e4ba5",
  1109 => x"fdfe49cb",
  1110 => x"c6c187ce",
  1111 => x"c1ffc087",
  1112 => x"cb49744a",
  1113 => x"eee1c191",
  1114 => x"c2797281",
  1115 => x"bf97deec",
  1116 => x"7487d802",
  1117 => x"c191de49",
  1118 => x"d9f1c284",
  1119 => x"c283714b",
  1120 => x"dd4adeec",
  1121 => x"dffcfe49",
  1122 => x"7487d887",
  1123 => x"c293de4b",
  1124 => x"cb83d9f1",
  1125 => x"51c049a3",
  1126 => x"6e7384c1",
  1127 => x"fe49cb4a",
  1128 => x"c487c5fc",
  1129 => x"80c14866",
  1130 => x"c758a6c8",
  1131 => x"c5c003ac",
  1132 => x"fc056e87",
  1133 => x"487487e0",
  1134 => x"fcf78ef4",
  1135 => x"1e731e87",
  1136 => x"cb494b71",
  1137 => x"eee1c191",
  1138 => x"4aa1c881",
  1139 => x"48d2e2c2",
  1140 => x"a1c95012",
  1141 => x"fcfdc04a",
  1142 => x"ca501248",
  1143 => x"d8f1c281",
  1144 => x"c2501148",
  1145 => x"bf97d8f1",
  1146 => x"49c01e49",
  1147 => x"87d3dac1",
  1148 => x"48c0f1c2",
  1149 => x"49c178de",
  1150 => x"2687cad6",
  1151 => x"1e87fef6",
  1152 => x"cb494a71",
  1153 => x"eee1c191",
  1154 => x"1181c881",
  1155 => x"c4f1c248",
  1156 => x"c4f1c258",
  1157 => x"c178c048",
  1158 => x"87e9d549",
  1159 => x"c01e4f26",
  1160 => x"e8c6c149",
  1161 => x"1e4f2687",
  1162 => x"d2029971",
  1163 => x"c3e3c187",
  1164 => x"f750c048",
  1165 => x"ffc7c180",
  1166 => x"e7e1c140",
  1167 => x"c187ce78",
  1168 => x"c148ffe2",
  1169 => x"fc78e0e1",
  1170 => x"dec8c180",
  1171 => x"0e4f2678",
  1172 => x"0e5c5b5e",
  1173 => x"cb4a4c71",
  1174 => x"eee1c192",
  1175 => x"49a2c882",
  1176 => x"974ba2c9",
  1177 => x"971e4b6b",
  1178 => x"ca1e4969",
  1179 => x"c0491282",
  1180 => x"c087c9e7",
  1181 => x"87cdd449",
  1182 => x"c3c14974",
  1183 => x"8ef887ea",
  1184 => x"1e87f8f4",
  1185 => x"4b711e73",
  1186 => x"87c3ff49",
  1187 => x"fefe4973",
  1188 => x"87e9f487",
  1189 => x"711e731e",
  1190 => x"4aa3c64b",
  1191 => x"c187db02",
  1192 => x"87d6028a",
  1193 => x"dac1028a",
  1194 => x"c0028a87",
  1195 => x"028a87fc",
  1196 => x"8a87e1c0",
  1197 => x"c187cb02",
  1198 => x"49c787db",
  1199 => x"c187c0fd",
  1200 => x"f1c287de",
  1201 => x"c102bfc4",
  1202 => x"c14887cb",
  1203 => x"c8f1c288",
  1204 => x"87c1c158",
  1205 => x"bfc8f1c2",
  1206 => x"87f9c002",
  1207 => x"bfc4f1c2",
  1208 => x"c280c148",
  1209 => x"c058c8f1",
  1210 => x"f1c287eb",
  1211 => x"c649bfc4",
  1212 => x"c8f1c289",
  1213 => x"a9b7c059",
  1214 => x"c287da03",
  1215 => x"c048c4f1",
  1216 => x"c287d278",
  1217 => x"02bfc8f1",
  1218 => x"f1c287cb",
  1219 => x"c648bfc4",
  1220 => x"c8f1c280",
  1221 => x"d149c058",
  1222 => x"497387eb",
  1223 => x"87c8c1c1",
  1224 => x"1e87daf2",
  1225 => x"4b711e73",
  1226 => x"48c0f1c2",
  1227 => x"49c078dd",
  1228 => x"7387d2d1",
  1229 => x"efc0c149",
  1230 => x"87c1f287",
  1231 => x"5c5b5e0e",
  1232 => x"cc4c710e",
  1233 => x"4b741e66",
  1234 => x"e1c193cb",
  1235 => x"a3c483ee",
  1236 => x"fe496a4a",
  1237 => x"c187e1f5",
  1238 => x"c87bfdc6",
  1239 => x"66d449a3",
  1240 => x"49a3c951",
  1241 => x"ca5166d8",
  1242 => x"66dc49a3",
  1243 => x"caf12651",
  1244 => x"5b5e0e87",
  1245 => x"ff0e5d5c",
  1246 => x"a6dc86cc",
  1247 => x"48a6c859",
  1248 => x"80c478c0",
  1249 => x"7866c8c1",
  1250 => x"78c180c4",
  1251 => x"78c180c4",
  1252 => x"48c8f1c2",
  1253 => x"f1c278c1",
  1254 => x"de48bfc0",
  1255 => x"87cb05a8",
  1256 => x"7087ccf3",
  1257 => x"59a6cc49",
  1258 => x"e787d6ce",
  1259 => x"c4e887d2",
  1260 => x"87ece687",
  1261 => x"fbc04c70",
  1262 => x"d8c102ac",
  1263 => x"0566d887",
  1264 => x"c087cac1",
  1265 => x"1ec11e1e",
  1266 => x"1ee1e3c1",
  1267 => x"ebfd49c0",
  1268 => x"c086d087",
  1269 => x"d902acfb",
  1270 => x"66c4c187",
  1271 => x"6a82c44a",
  1272 => x"7481c749",
  1273 => x"d81ec151",
  1274 => x"c8496a1e",
  1275 => x"87d9e781",
  1276 => x"c8c186c8",
  1277 => x"a8c04866",
  1278 => x"c887c701",
  1279 => x"78c148a6",
  1280 => x"c8c187ce",
  1281 => x"88c14866",
  1282 => x"c358a6d0",
  1283 => x"87e5e687",
  1284 => x"c248a6d0",
  1285 => x"029c7478",
  1286 => x"c887e2cc",
  1287 => x"ccc14866",
  1288 => x"cc03a866",
  1289 => x"a6dc87d7",
  1290 => x"e478c048",
  1291 => x"4c7087f2",
  1292 => x"dd4866d8",
  1293 => x"87c605a8",
  1294 => x"d848a6dc",
  1295 => x"d0c17866",
  1296 => x"e8c005ac",
  1297 => x"87d8e487",
  1298 => x"7087d5e4",
  1299 => x"acecc04c",
  1300 => x"e587c505",
  1301 => x"4c7087df",
  1302 => x"05acd0c1",
  1303 => x"66d487c8",
  1304 => x"d880c148",
  1305 => x"d0c158a6",
  1306 => x"d8ff02ac",
  1307 => x"a6e0c087",
  1308 => x"7866d848",
  1309 => x"c04866dc",
  1310 => x"05a866e0",
  1311 => x"c487d0ca",
  1312 => x"f0c048a6",
  1313 => x"80e0c078",
  1314 => x"c47866d0",
  1315 => x"c478c080",
  1316 => x"7478c080",
  1317 => x"8dfbc04d",
  1318 => x"87ccc902",
  1319 => x"db028dc9",
  1320 => x"028dc287",
  1321 => x"c987cdc1",
  1322 => x"d1c4028d",
  1323 => x"028dc487",
  1324 => x"c187cec1",
  1325 => x"c5c4028d",
  1326 => x"87e6c887",
  1327 => x"cb4966c8",
  1328 => x"66c4c191",
  1329 => x"4aa1c481",
  1330 => x"1e717e6a",
  1331 => x"48f8ddc1",
  1332 => x"cc4966c4",
  1333 => x"41204aa1",
  1334 => x"ff05aa71",
  1335 => x"511087f8",
  1336 => x"ccc14926",
  1337 => x"cce379e3",
  1338 => x"c04c7087",
  1339 => x"c148a6ec",
  1340 => x"87f4c778",
  1341 => x"c048a6c4",
  1342 => x"4866d078",
  1343 => x"a6d480c1",
  1344 => x"87dce158",
  1345 => x"ecc04c70",
  1346 => x"87d402ac",
  1347 => x"c00266c4",
  1348 => x"a6c887c5",
  1349 => x"7487c95c",
  1350 => x"88f0c048",
  1351 => x"58a6e8c0",
  1352 => x"02acecc0",
  1353 => x"f7e087cc",
  1354 => x"c04c7087",
  1355 => x"ff05acec",
  1356 => x"66c487f4",
  1357 => x"4966d81e",
  1358 => x"66ecc01e",
  1359 => x"e1e3c11e",
  1360 => x"4966d81e",
  1361 => x"c087f5f7",
  1362 => x"c01eca1e",
  1363 => x"cb4966e0",
  1364 => x"66dcc191",
  1365 => x"48a6d881",
  1366 => x"d878a1c4",
  1367 => x"e149bf66",
  1368 => x"86d887e7",
  1369 => x"06a8b7c0",
  1370 => x"c187cac1",
  1371 => x"c81ede1e",
  1372 => x"e149bf66",
  1373 => x"86c887d3",
  1374 => x"c0484970",
  1375 => x"e8c08808",
  1376 => x"b7c058a6",
  1377 => x"ecc006a8",
  1378 => x"66e4c087",
  1379 => x"a8b7dd48",
  1380 => x"87e1c003",
  1381 => x"c049bf6e",
  1382 => x"c08166e4",
  1383 => x"e4c051e0",
  1384 => x"81c14966",
  1385 => x"c281bf6e",
  1386 => x"e4c051c1",
  1387 => x"81c24966",
  1388 => x"c081bf6e",
  1389 => x"a6ecc051",
  1390 => x"c478c148",
  1391 => x"f7e187ea",
  1392 => x"a6e8c087",
  1393 => x"87f0e158",
  1394 => x"58a6f0c0",
  1395 => x"05a8ecc0",
  1396 => x"a687c9c0",
  1397 => x"66e4c048",
  1398 => x"87c4c078",
  1399 => x"87c0deff",
  1400 => x"cb4966c8",
  1401 => x"66c4c191",
  1402 => x"c8807148",
  1403 => x"66c458a6",
  1404 => x"c482c84a",
  1405 => x"81ca4966",
  1406 => x"5166e4c0",
  1407 => x"4966ecc0",
  1408 => x"e4c081c1",
  1409 => x"48c18966",
  1410 => x"49703071",
  1411 => x"977189c1",
  1412 => x"f5f4c27a",
  1413 => x"e4c049bf",
  1414 => x"6a972966",
  1415 => x"9871484a",
  1416 => x"58a6f4c0",
  1417 => x"c44966c4",
  1418 => x"c07e6981",
  1419 => x"dc4866e0",
  1420 => x"c002a866",
  1421 => x"a6dc87c8",
  1422 => x"c078c048",
  1423 => x"a6dc87c5",
  1424 => x"dc78c148",
  1425 => x"e0c01e66",
  1426 => x"4966c81e",
  1427 => x"87f9ddff",
  1428 => x"4c7086c8",
  1429 => x"06acb7c0",
  1430 => x"6e87d6c1",
  1431 => x"70807448",
  1432 => x"49e0c07e",
  1433 => x"4b6e8974",
  1434 => x"4af5ddc1",
  1435 => x"f7e8fe71",
  1436 => x"c2486e87",
  1437 => x"c07e7080",
  1438 => x"c14866e8",
  1439 => x"a6ecc080",
  1440 => x"66f0c058",
  1441 => x"7081c149",
  1442 => x"c5c002a9",
  1443 => x"c04dc087",
  1444 => x"4dc187c2",
  1445 => x"a4c21e75",
  1446 => x"48e0c049",
  1447 => x"49708871",
  1448 => x"4966c81e",
  1449 => x"87e1dcff",
  1450 => x"b7c086c8",
  1451 => x"c6ff01a8",
  1452 => x"66e8c087",
  1453 => x"87d3c002",
  1454 => x"c94966c4",
  1455 => x"66e8c081",
  1456 => x"4866c451",
  1457 => x"78cfc9c1",
  1458 => x"c487cec0",
  1459 => x"81c94966",
  1460 => x"66c451c2",
  1461 => x"c3cac148",
  1462 => x"a6ecc078",
  1463 => x"c078c148",
  1464 => x"dbff87c6",
  1465 => x"4c7087cf",
  1466 => x"0266ecc0",
  1467 => x"c887f5c0",
  1468 => x"66cc4866",
  1469 => x"cbc004a8",
  1470 => x"4866c887",
  1471 => x"a6cc80c1",
  1472 => x"87e0c058",
  1473 => x"c14866cc",
  1474 => x"58a6d088",
  1475 => x"c187d5c0",
  1476 => x"c005acc6",
  1477 => x"66d087c8",
  1478 => x"d480c148",
  1479 => x"daff58a6",
  1480 => x"4c7087d3",
  1481 => x"c14866d4",
  1482 => x"58a6d880",
  1483 => x"c0029c74",
  1484 => x"66c887cb",
  1485 => x"66ccc148",
  1486 => x"e9f304a8",
  1487 => x"ebd9ff87",
  1488 => x"4866c887",
  1489 => x"c003a8c7",
  1490 => x"f1c287e5",
  1491 => x"78c048c8",
  1492 => x"cb4966c8",
  1493 => x"66c4c191",
  1494 => x"4aa1c481",
  1495 => x"52c04a6a",
  1496 => x"4866c879",
  1497 => x"a6cc80c1",
  1498 => x"04a8c758",
  1499 => x"ff87dbff",
  1500 => x"c4e18ecc",
  1501 => x"00203a87",
  1502 => x"20504944",
  1503 => x"74697753",
  1504 => x"73656863",
  1505 => x"1e731e00",
  1506 => x"029b4b71",
  1507 => x"f1c287c6",
  1508 => x"78c048c4",
  1509 => x"f1c21ec7",
  1510 => x"1e49bfc4",
  1511 => x"1eeee1c1",
  1512 => x"bfc0f1c2",
  1513 => x"87c9ef49",
  1514 => x"f1c286cc",
  1515 => x"e949bfc0",
  1516 => x"9b7387f5",
  1517 => x"c187c802",
  1518 => x"c049eee1",
  1519 => x"ff87fbef",
  1520 => x"1e87fadf",
  1521 => x"48d2e2c2",
  1522 => x"e3c150c0",
  1523 => x"c049bfd1",
  1524 => x"c087c7fe",
  1525 => x"1e4f2648",
  1526 => x"c187e5c7",
  1527 => x"87e5fe49",
  1528 => x"87ceebfe",
  1529 => x"cd029870",
  1530 => x"e9f2fe87",
  1531 => x"02987087",
  1532 => x"4ac187c4",
  1533 => x"4ac087c2",
  1534 => x"ce059a72",
  1535 => x"c11ec087",
  1536 => x"c049ebe0",
  1537 => x"c487d1fb",
  1538 => x"c187fe86",
  1539 => x"c087edc2",
  1540 => x"f6e0c11e",
  1541 => x"fffac049",
  1542 => x"fe1ec087",
  1543 => x"497087e5",
  1544 => x"87f4fac0",
  1545 => x"f887d8c3",
  1546 => x"534f268e",
  1547 => x"61662044",
  1548 => x"64656c69",
  1549 => x"6f42002e",
  1550 => x"6e69746f",
  1551 => x"2e2e2e67",
  1552 => x"f2c01e00",
  1553 => x"87fa87d5",
  1554 => x"c21e4f26",
  1555 => x"c048c4f1",
  1556 => x"c0f1c278",
  1557 => x"fd78c048",
  1558 => x"87e587fd",
  1559 => x"4f2648c0",
  1560 => x"78452080",
  1561 => x"80007469",
  1562 => x"63614220",
  1563 => x"11ff006b",
  1564 => x"2c590000",
  1565 => x"00000000",
  1566 => x"0011ff00",
  1567 => x"002c7700",
  1568 => x"00000000",
  1569 => x"000011ff",
  1570 => x"00002c95",
  1571 => x"ff000000",
  1572 => x"b3000011",
  1573 => x"0000002c",
  1574 => x"11ff0000",
  1575 => x"2cd10000",
  1576 => x"00000000",
  1577 => x"0011ff00",
  1578 => x"002cef00",
  1579 => x"00000000",
  1580 => x"000011ff",
  1581 => x"00002d0d",
  1582 => x"ff000000",
  1583 => x"00000011",
  1584 => x"00000000",
  1585 => x"12940000",
  1586 => x"00000000",
  1587 => x"00000000",
  1588 => x"0018d500",
  1589 => x"4f4f4200",
  1590 => x"20202054",
  1591 => x"4d4f5220",
  1592 => x"616f4c00",
  1593 => x"2e2a2064",
  1594 => x"f0fe1e00",
  1595 => x"cd78c048",
  1596 => x"26097909",
  1597 => x"fe1e1e4f",
  1598 => x"487ebff0",
  1599 => x"1e4f2626",
  1600 => x"c148f0fe",
  1601 => x"1e4f2678",
  1602 => x"c048f0fe",
  1603 => x"1e4f2678",
  1604 => x"52c04a71",
  1605 => x"0e4f2652",
  1606 => x"5d5c5b5e",
  1607 => x"7186f40e",
  1608 => x"7e6d974d",
  1609 => x"974ca5c1",
  1610 => x"a6c8486c",
  1611 => x"c4486e58",
  1612 => x"c505a866",
  1613 => x"c048ff87",
  1614 => x"caff87e6",
  1615 => x"49a5c287",
  1616 => x"714b6c97",
  1617 => x"6b974ba3",
  1618 => x"7e6c974b",
  1619 => x"80c1486e",
  1620 => x"c758a6c8",
  1621 => x"58a6cc98",
  1622 => x"fe7c9770",
  1623 => x"487387e1",
  1624 => x"4d268ef4",
  1625 => x"4b264c26",
  1626 => x"5e0e4f26",
  1627 => x"f40e5c5b",
  1628 => x"d84c7186",
  1629 => x"ffc34a66",
  1630 => x"4ba4c29a",
  1631 => x"73496c97",
  1632 => x"517249a1",
  1633 => x"6e7e6c97",
  1634 => x"c880c148",
  1635 => x"98c758a6",
  1636 => x"7058a6cc",
  1637 => x"ff8ef454",
  1638 => x"1e1e87ca",
  1639 => x"e087e8fd",
  1640 => x"c0494abf",
  1641 => x"0299c0e0",
  1642 => x"1e7287cb",
  1643 => x"49ebf4c2",
  1644 => x"c487f7fe",
  1645 => x"87fdfc86",
  1646 => x"c2fd7e70",
  1647 => x"4f262687",
  1648 => x"ebf4c21e",
  1649 => x"87c7fd49",
  1650 => x"49dae6c1",
  1651 => x"c587dafc",
  1652 => x"4f2687d9",
  1653 => x"5c5b5e0e",
  1654 => x"f5c20e5d",
  1655 => x"c14abffe",
  1656 => x"49bfe8e8",
  1657 => x"71bc724c",
  1658 => x"87dbfc4d",
  1659 => x"49744bc0",
  1660 => x"d50299d0",
  1661 => x"d0497587",
  1662 => x"c01e7199",
  1663 => x"faeec11e",
  1664 => x"1282734a",
  1665 => x"87e4c049",
  1666 => x"2cc186c8",
  1667 => x"abc8832d",
  1668 => x"87daff04",
  1669 => x"c187e8fb",
  1670 => x"c248e8e8",
  1671 => x"78bffef5",
  1672 => x"4c264d26",
  1673 => x"4f264b26",
  1674 => x"00000000",
  1675 => x"48d0ff1e",
  1676 => x"ff78e1c8",
  1677 => x"78c548d4",
  1678 => x"c30266c4",
  1679 => x"78e0c387",
  1680 => x"c60266c8",
  1681 => x"48d4ff87",
  1682 => x"ff78f0c3",
  1683 => x"787148d4",
  1684 => x"c848d0ff",
  1685 => x"e0c078e1",
  1686 => x"0e4f2678",
  1687 => x"0e5c5b5e",
  1688 => x"f4c24c71",
  1689 => x"eefa49eb",
  1690 => x"c04a7087",
  1691 => x"c204aab7",
  1692 => x"e0c387e3",
  1693 => x"87c905aa",
  1694 => x"48deecc1",
  1695 => x"d4c278c1",
  1696 => x"aaf0c387",
  1697 => x"c187c905",
  1698 => x"c148daec",
  1699 => x"87f5c178",
  1700 => x"bfdeecc1",
  1701 => x"7287c702",
  1702 => x"b3c0c24b",
  1703 => x"4b7287c2",
  1704 => x"d1059c74",
  1705 => x"daecc187",
  1706 => x"ecc11ebf",
  1707 => x"721ebfde",
  1708 => x"87f8fd49",
  1709 => x"ecc186c8",
  1710 => x"c002bfda",
  1711 => x"497387e0",
  1712 => x"9129b7c4",
  1713 => x"81faedc1",
  1714 => x"9acf4a73",
  1715 => x"48c192c2",
  1716 => x"4a703072",
  1717 => x"4872baff",
  1718 => x"79709869",
  1719 => x"497387db",
  1720 => x"9129b7c4",
  1721 => x"81faedc1",
  1722 => x"9acf4a73",
  1723 => x"48c392c2",
  1724 => x"4a703072",
  1725 => x"70b06948",
  1726 => x"deecc179",
  1727 => x"c178c048",
  1728 => x"c048daec",
  1729 => x"ebf4c278",
  1730 => x"87cbf849",
  1731 => x"b7c04a70",
  1732 => x"ddfd03aa",
  1733 => x"fc48c087",
  1734 => x"000087c8",
  1735 => x"00000000",
  1736 => x"711e0000",
  1737 => x"f2fc494a",
  1738 => x"1e4f2687",
  1739 => x"49724ac0",
  1740 => x"edc191c4",
  1741 => x"79c081fa",
  1742 => x"b7d082c1",
  1743 => x"87ee04aa",
  1744 => x"5e0e4f26",
  1745 => x"0e5d5c5b",
  1746 => x"faf64d71",
  1747 => x"c44a7587",
  1748 => x"c1922ab7",
  1749 => x"7582faed",
  1750 => x"c29ccf4c",
  1751 => x"4b496a94",
  1752 => x"9bc32b74",
  1753 => x"307448c2",
  1754 => x"bcff4c70",
  1755 => x"98714874",
  1756 => x"caf67a70",
  1757 => x"fa487387",
  1758 => x"000087e6",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"1e160000",
  1775 => x"362e2526",
  1776 => x"ff1e3e3d",
  1777 => x"e1c848d0",
  1778 => x"ff487178",
  1779 => x"c47808d4",
  1780 => x"d4ff4866",
  1781 => x"4f267808",
  1782 => x"c44a711e",
  1783 => x"721e4966",
  1784 => x"87deff49",
  1785 => x"c048d0ff",
  1786 => x"262678e0",
  1787 => x"4a711e4f",
  1788 => x"c11e66c4",
  1789 => x"ff49a2e0",
  1790 => x"66c887c8",
  1791 => x"29b7c849",
  1792 => x"7148d4ff",
  1793 => x"48d0ff78",
  1794 => x"2678e0c0",
  1795 => x"ff1e4f26",
  1796 => x"ffc34ad4",
  1797 => x"48d0ff7a",
  1798 => x"de78e1c8",
  1799 => x"f5f4c27a",
  1800 => x"48497abf",
  1801 => x"7a7028c8",
  1802 => x"28d04871",
  1803 => x"48717a70",
  1804 => x"7a7028d8",
  1805 => x"c048d0ff",
  1806 => x"4f2678e0",
  1807 => x"5c5b5e0e",
  1808 => x"4c710e5d",
  1809 => x"bff5f4c2",
  1810 => x"2b744b4d",
  1811 => x"c19b66d0",
  1812 => x"ab66d483",
  1813 => x"c087c204",
  1814 => x"d04a744b",
  1815 => x"31724966",
  1816 => x"9975b9ff",
  1817 => x"30724873",
  1818 => x"71484a70",
  1819 => x"f9f4c2b0",
  1820 => x"87dafe58",
  1821 => x"4c264d26",
  1822 => x"4f264b26",
  1823 => x"5c5b5e0e",
  1824 => x"711e0e5d",
  1825 => x"f9f4c24c",
  1826 => x"c04ac04b",
  1827 => x"d0fe49f4",
  1828 => x"1e7487f3",
  1829 => x"49f9f4c2",
  1830 => x"87c6edfe",
  1831 => x"987086c4",
  1832 => x"87eac002",
  1833 => x"4da61ec4",
  1834 => x"f9f4c21e",
  1835 => x"f7f2fe49",
  1836 => x"7086c887",
  1837 => x"87d60298",
  1838 => x"f4c14a75",
  1839 => x"4bc449c4",
  1840 => x"87e6cefe",
  1841 => x"ca029870",
  1842 => x"c048c087",
  1843 => x"48c087ed",
  1844 => x"c087e8c0",
  1845 => x"c4c187f3",
  1846 => x"02987087",
  1847 => x"fcc087c8",
  1848 => x"05987087",
  1849 => x"f5c287f8",
  1850 => x"cc02bfd9",
  1851 => x"f5f4c287",
  1852 => x"d9f5c248",
  1853 => x"d5fc78bf",
  1854 => x"2648c187",
  1855 => x"4c264d26",
  1856 => x"4f264b26",
  1857 => x"4352415b",
  1858 => x"1ec01e00",
  1859 => x"49f9f4c2",
  1860 => x"87edeffe",
  1861 => x"48d1f5c2",
  1862 => x"262678c0",
  1863 => x"5b5e0e4f",
  1864 => x"f40e5d5c",
  1865 => x"48a6c486",
  1866 => x"f5c278c0",
  1867 => x"c348bfd1",
  1868 => x"d103a8b7",
  1869 => x"d1f5c287",
  1870 => x"80c148bf",
  1871 => x"58d5f5c2",
  1872 => x"c648fbc0",
  1873 => x"f4c287e2",
  1874 => x"f4fe49f9",
  1875 => x"4c7087ee",
  1876 => x"bfd1f5c2",
  1877 => x"028ac34a",
  1878 => x"8ac187d8",
  1879 => x"87cbc502",
  1880 => x"f6c2028a",
  1881 => x"c1028a87",
  1882 => x"028a87cd",
  1883 => x"c587e2c3",
  1884 => x"4dc087e1",
  1885 => x"92c44a75",
  1886 => x"82c6fcc1",
  1887 => x"48cdf5c2",
  1888 => x"7e708075",
  1889 => x"4bbf976e",
  1890 => x"486e4b49",
  1891 => x"6a50a3c1",
  1892 => x"cc481181",
  1893 => x"ac7058a6",
  1894 => x"6e87c402",
  1895 => x"c850c048",
  1896 => x"87c70566",
  1897 => x"48d1f5c2",
  1898 => x"c178a5c4",
  1899 => x"adb7c485",
  1900 => x"87c0ff04",
  1901 => x"c287dcc4",
  1902 => x"48bfddf5",
  1903 => x"01a8b7c8",
  1904 => x"acca87d1",
  1905 => x"cd87cc02",
  1906 => x"87c702ac",
  1907 => x"03acb7c0",
  1908 => x"c287f3c0",
  1909 => x"4bbfddf5",
  1910 => x"03abb7c8",
  1911 => x"f5c287d2",
  1912 => x"817349e1",
  1913 => x"c151e0c0",
  1914 => x"abb7c883",
  1915 => x"87eeff04",
  1916 => x"48e9f5c2",
  1917 => x"c150d2c1",
  1918 => x"cdc150cf",
  1919 => x"e450c050",
  1920 => x"c378c380",
  1921 => x"f5c287cd",
  1922 => x"4849bfdd",
  1923 => x"f5c280c1",
  1924 => x"c44858e1",
  1925 => x"517481a0",
  1926 => x"c087f8c2",
  1927 => x"04acb7f0",
  1928 => x"f9c087da",
  1929 => x"d301acb7",
  1930 => x"d5f5c287",
  1931 => x"91ca49bf",
  1932 => x"f0c04a74",
  1933 => x"d5f5c28a",
  1934 => x"78a17248",
  1935 => x"c002acca",
  1936 => x"accd87c6",
  1937 => x"87cbc205",
  1938 => x"48d1f5c2",
  1939 => x"c2c278c3",
  1940 => x"b7f0c087",
  1941 => x"87db04ac",
  1942 => x"acb7f9c0",
  1943 => x"87d3c001",
  1944 => x"bfd9f5c2",
  1945 => x"7491d049",
  1946 => x"8af0c04a",
  1947 => x"48d9f5c2",
  1948 => x"c178a172",
  1949 => x"04acb7c1",
  1950 => x"c187dbc0",
  1951 => x"01acb7c6",
  1952 => x"c287d3c0",
  1953 => x"49bfd9f5",
  1954 => x"4a7491d0",
  1955 => x"c28af7c0",
  1956 => x"7248d9f5",
  1957 => x"acca78a1",
  1958 => x"87c6c002",
  1959 => x"c005accd",
  1960 => x"f5c287f1",
  1961 => x"78c348d1",
  1962 => x"c087e8c0",
  1963 => x"c005ace2",
  1964 => x"a6c487c9",
  1965 => x"78fbc048",
  1966 => x"ca87d8c0",
  1967 => x"c6c002ac",
  1968 => x"05accd87",
  1969 => x"c287c9c0",
  1970 => x"c348d1f5",
  1971 => x"87c3c078",
  1972 => x"c05ca6c8",
  1973 => x"c003acb7",
  1974 => x"c04887c4",
  1975 => x"66c487ca",
  1976 => x"87c6f902",
  1977 => x"99ffc348",
  1978 => x"cff88ef4",
  1979 => x"4e4f4387",
  1980 => x"4d003d46",
  1981 => x"4e00444f",
  1982 => x"00454d41",
  1983 => x"41464544",
  1984 => x"3d544c55",
  1985 => x"1eed0030",
  1986 => x"1ef30000",
  1987 => x"1ef70000",
  1988 => x"1efc0000",
  1989 => x"ff1e0000",
  1990 => x"c9c848d0",
  1991 => x"ff487178",
  1992 => x"267808d4",
  1993 => x"4a711e4f",
  1994 => x"ff87eb49",
  1995 => x"78c848d0",
  1996 => x"731e4f26",
  1997 => x"c24b711e",
  1998 => x"02bff9f5",
  1999 => x"ebc287c3",
  2000 => x"48d0ff87",
  2001 => x"7378c9c8",
  2002 => x"b1e0c049",
  2003 => x"7148d4ff",
  2004 => x"edf5c278",
  2005 => x"c878c048",
  2006 => x"87c50266",
  2007 => x"c249ffc3",
  2008 => x"c249c087",
  2009 => x"cc59f5f5",
  2010 => x"87c60266",
  2011 => x"4ad5d5c5",
  2012 => x"ffcf87c4",
  2013 => x"f5c24aff",
  2014 => x"f5c25af9",
  2015 => x"78c148f9",
  2016 => x"4d2687c4",
  2017 => x"4b264c26",
  2018 => x"5e0e4f26",
  2019 => x"0e5d5c5b",
  2020 => x"f5c24a71",
  2021 => x"724cbff5",
  2022 => x"87cb029a",
  2023 => x"c191c849",
  2024 => x"714be8fc",
  2025 => x"c287c483",
  2026 => x"c04be8c0",
  2027 => x"7449134d",
  2028 => x"f1f5c299",
  2029 => x"d4ffb9bf",
  2030 => x"c1787148",
  2031 => x"c8852cb7",
  2032 => x"e804adb7",
  2033 => x"edf5c287",
  2034 => x"80c848bf",
  2035 => x"58f1f5c2",
  2036 => x"1e87effe",
  2037 => x"4b711e73",
  2038 => x"029a4a13",
  2039 => x"497287cb",
  2040 => x"1387e7fe",
  2041 => x"f5059a4a",
  2042 => x"87dafe87",
  2043 => x"edf5c21e",
  2044 => x"f5c249bf",
  2045 => x"a1c148ed",
  2046 => x"b7c0c478",
  2047 => x"87db03a9",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
